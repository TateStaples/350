

module wallaceTreeMultiplier(
    data_operandA, data_operandB, 
    clock, 
    data_result, data_exception, data_resultRDY);

    input [31:0] data_operandA, data_operandB;
    input clock;

    output [63:0] data_result;
    output data_exception, data_resultRDY;

    assign data_resultRDY = 1'b1;

wire [31:0] partialProduct_0, partialProduct_1, partialProduct_2, partialProduct_3, partialProduct_4, partialProduct_5, partialProduct_6, partialProduct_7, partialProduct_8, partialProduct_9, partialProduct_10, partialProduct_11, partialProduct_12, partialProduct_13, partialProduct_14, partialProduct_15, partialProduct_16, partialProduct_17, partialProduct_18, partialProduct_19, partialProduct_20, partialProduct_21, partialProduct_22, partialProduct_23, partialProduct_24, partialProduct_25, partialProduct_26, partialProduct_27, partialProduct_28, partialProduct_29, partialProduct_30, partialProduct_31;
assign partialProduct_0 = data_operandA & {32{data_operandB[0]}};
assign partialProduct_1 = data_operandA & {32{data_operandB[1]}};
assign partialProduct_2 = data_operandA & {32{data_operandB[2]}};
assign partialProduct_3 = data_operandA & {32{data_operandB[3]}};
assign partialProduct_4 = data_operandA & {32{data_operandB[4]}};
assign partialProduct_5 = data_operandA & {32{data_operandB[5]}};
assign partialProduct_6 = data_operandA & {32{data_operandB[6]}};
assign partialProduct_7 = data_operandA & {32{data_operandB[7]}};
assign partialProduct_8 = data_operandA & {32{data_operandB[8]}};
assign partialProduct_9 = data_operandA & {32{data_operandB[9]}};
assign partialProduct_10 = data_operandA & {32{data_operandB[10]}};
assign partialProduct_11 = data_operandA & {32{data_operandB[11]}};
assign partialProduct_12 = data_operandA & {32{data_operandB[12]}};
assign partialProduct_13 = data_operandA & {32{data_operandB[13]}};
assign partialProduct_14 = data_operandA & {32{data_operandB[14]}};
assign partialProduct_15 = data_operandA & {32{data_operandB[15]}};
assign partialProduct_16 = data_operandA & {32{data_operandB[16]}};
assign partialProduct_17 = data_operandA & {32{data_operandB[17]}};
assign partialProduct_18 = data_operandA & {32{data_operandB[18]}};
assign partialProduct_19 = data_operandA & {32{data_operandB[19]}};
assign partialProduct_20 = data_operandA & {32{data_operandB[20]}};
assign partialProduct_21 = data_operandA & {32{data_operandB[21]}};
assign partialProduct_22 = data_operandA & {32{data_operandB[22]}};
assign partialProduct_23 = data_operandA & {32{data_operandB[23]}};
assign partialProduct_24 = data_operandA & {32{data_operandB[24]}};
assign partialProduct_25 = data_operandA & {32{data_operandB[25]}};
assign partialProduct_26 = data_operandA & {32{data_operandB[26]}};
assign partialProduct_27 = data_operandA & {32{data_operandB[27]}};
assign partialProduct_28 = data_operandA & {32{data_operandB[28]}};
assign partialProduct_29 = data_operandA & {32{data_operandB[29]}};
assign partialProduct_30 = data_operandA & {32{data_operandB[30]}};
assign partialProduct_31 = data_operandA & {32{data_operandB[31]}};
wire wire_0, wire_1;
assign wire_0 = partialProduct_0[1] ^ partialProduct_1[0];
assign wire_1 = partialProduct_0[1] & partialProduct_1[0];
wire wire_2, wire_3;
bit_adder add0(.S(wire_2), .Cout(wire_3),  .A(partialProduct_0[2]), .B(partialProduct_1[1]), .Cin(partialProduct_2[0]));
wire wire_4, wire_5;
bit_adder add1(.S(wire_4), .Cout(wire_5),  .A(partialProduct_0[3]), .B(partialProduct_1[2]), .Cin(partialProduct_2[1]));
wire wire_6, wire_7;
bit_adder add2(.S(wire_6), .Cout(wire_7),  .A(partialProduct_0[4]), .B(partialProduct_1[3]), .Cin(partialProduct_2[2]));
wire wire_8, wire_9;
bit_adder add3(.S(wire_8), .Cout(wire_9),  .A(partialProduct_0[5]), .B(partialProduct_1[4]), .Cin(partialProduct_2[3]));
wire wire_10, wire_11;
bit_adder add4(.S(wire_10), .Cout(wire_11),  .A(partialProduct_0[6]), .B(partialProduct_1[5]), .Cin(partialProduct_2[4]));
wire wire_12, wire_13;
bit_adder add5(.S(wire_12), .Cout(wire_13),  .A(partialProduct_0[7]), .B(partialProduct_1[6]), .Cin(partialProduct_2[5]));
wire wire_14, wire_15;
bit_adder add6(.S(wire_14), .Cout(wire_15),  .A(partialProduct_0[8]), .B(partialProduct_1[7]), .Cin(partialProduct_2[6]));
wire wire_16, wire_17;
bit_adder add7(.S(wire_16), .Cout(wire_17),  .A(partialProduct_0[9]), .B(partialProduct_1[8]), .Cin(partialProduct_2[7]));
wire wire_18, wire_19;
bit_adder add8(.S(wire_18), .Cout(wire_19),  .A(partialProduct_0[10]), .B(partialProduct_1[9]), .Cin(partialProduct_2[8]));
wire wire_20, wire_21;
bit_adder add9(.S(wire_20), .Cout(wire_21),  .A(partialProduct_0[11]), .B(partialProduct_1[10]), .Cin(partialProduct_2[9]));
wire wire_22, wire_23;
bit_adder add10(.S(wire_22), .Cout(wire_23),  .A(partialProduct_0[12]), .B(partialProduct_1[11]), .Cin(partialProduct_2[10]));
wire wire_24, wire_25;
bit_adder add11(.S(wire_24), .Cout(wire_25),  .A(partialProduct_0[13]), .B(partialProduct_1[12]), .Cin(partialProduct_2[11]));
wire wire_26, wire_27;
bit_adder add12(.S(wire_26), .Cout(wire_27),  .A(partialProduct_0[14]), .B(partialProduct_1[13]), .Cin(partialProduct_2[12]));
wire wire_28, wire_29;
bit_adder add13(.S(wire_28), .Cout(wire_29),  .A(partialProduct_0[15]), .B(partialProduct_1[14]), .Cin(partialProduct_2[13]));
wire wire_30, wire_31;
bit_adder add14(.S(wire_30), .Cout(wire_31),  .A(partialProduct_0[16]), .B(partialProduct_1[15]), .Cin(partialProduct_2[14]));
wire wire_32, wire_33;
bit_adder add15(.S(wire_32), .Cout(wire_33),  .A(partialProduct_0[17]), .B(partialProduct_1[16]), .Cin(partialProduct_2[15]));
wire wire_34, wire_35;
bit_adder add16(.S(wire_34), .Cout(wire_35),  .A(partialProduct_0[18]), .B(partialProduct_1[17]), .Cin(partialProduct_2[16]));
wire wire_36, wire_37;
bit_adder add17(.S(wire_36), .Cout(wire_37),  .A(partialProduct_0[19]), .B(partialProduct_1[18]), .Cin(partialProduct_2[17]));
wire wire_38, wire_39;
bit_adder add18(.S(wire_38), .Cout(wire_39),  .A(partialProduct_0[20]), .B(partialProduct_1[19]), .Cin(partialProduct_2[18]));
wire wire_40, wire_41;
bit_adder add19(.S(wire_40), .Cout(wire_41),  .A(partialProduct_0[21]), .B(partialProduct_1[20]), .Cin(partialProduct_2[19]));
wire wire_42, wire_43;
bit_adder add20(.S(wire_42), .Cout(wire_43),  .A(partialProduct_0[22]), .B(partialProduct_1[21]), .Cin(partialProduct_2[20]));
wire wire_44, wire_45;
bit_adder add21(.S(wire_44), .Cout(wire_45),  .A(partialProduct_0[23]), .B(partialProduct_1[22]), .Cin(partialProduct_2[21]));
wire wire_46, wire_47;
bit_adder add22(.S(wire_46), .Cout(wire_47),  .A(partialProduct_0[24]), .B(partialProduct_1[23]), .Cin(partialProduct_2[22]));
wire wire_48, wire_49;
bit_adder add23(.S(wire_48), .Cout(wire_49),  .A(partialProduct_0[25]), .B(partialProduct_1[24]), .Cin(partialProduct_2[23]));
wire wire_50, wire_51;
bit_adder add24(.S(wire_50), .Cout(wire_51),  .A(partialProduct_0[26]), .B(partialProduct_1[25]), .Cin(partialProduct_2[24]));
wire wire_52, wire_53;
bit_adder add25(.S(wire_52), .Cout(wire_53),  .A(partialProduct_0[27]), .B(partialProduct_1[26]), .Cin(partialProduct_2[25]));
wire wire_54, wire_55;
bit_adder add26(.S(wire_54), .Cout(wire_55),  .A(partialProduct_0[28]), .B(partialProduct_1[27]), .Cin(partialProduct_2[26]));
wire wire_56, wire_57;
bit_adder add27(.S(wire_56), .Cout(wire_57),  .A(partialProduct_0[29]), .B(partialProduct_1[28]), .Cin(partialProduct_2[27]));
wire wire_58, wire_59;
bit_adder add28(.S(wire_58), .Cout(wire_59),  .A(partialProduct_0[30]), .B(partialProduct_1[29]), .Cin(partialProduct_2[28]));
wire wire_60, wire_61;
bit_adder add29(.S(wire_60), .Cout(wire_61),  .A(partialProduct_0[31]), .B(partialProduct_1[30]), .Cin(partialProduct_2[29]));
wire wire_62, wire_63;
assign wire_62 = partialProduct_1[31] ^ partialProduct_2[30];
assign wire_63 = partialProduct_1[31] & partialProduct_2[30];
wire wire_64, wire_65;
assign wire_64 = partialProduct_3[1] ^ partialProduct_4[0];
assign wire_65 = partialProduct_3[1] & partialProduct_4[0];
wire wire_66, wire_67;
bit_adder add30(.S(wire_66), .Cout(wire_67),  .A(partialProduct_3[2]), .B(partialProduct_4[1]), .Cin(partialProduct_5[0]));
wire wire_68, wire_69;
bit_adder add31(.S(wire_68), .Cout(wire_69),  .A(partialProduct_3[3]), .B(partialProduct_4[2]), .Cin(partialProduct_5[1]));
wire wire_70, wire_71;
bit_adder add32(.S(wire_70), .Cout(wire_71),  .A(partialProduct_3[4]), .B(partialProduct_4[3]), .Cin(partialProduct_5[2]));
wire wire_72, wire_73;
bit_adder add33(.S(wire_72), .Cout(wire_73),  .A(partialProduct_3[5]), .B(partialProduct_4[4]), .Cin(partialProduct_5[3]));
wire wire_74, wire_75;
bit_adder add34(.S(wire_74), .Cout(wire_75),  .A(partialProduct_3[6]), .B(partialProduct_4[5]), .Cin(partialProduct_5[4]));
wire wire_76, wire_77;
bit_adder add35(.S(wire_76), .Cout(wire_77),  .A(partialProduct_3[7]), .B(partialProduct_4[6]), .Cin(partialProduct_5[5]));
wire wire_78, wire_79;
bit_adder add36(.S(wire_78), .Cout(wire_79),  .A(partialProduct_3[8]), .B(partialProduct_4[7]), .Cin(partialProduct_5[6]));
wire wire_80, wire_81;
bit_adder add37(.S(wire_80), .Cout(wire_81),  .A(partialProduct_3[9]), .B(partialProduct_4[8]), .Cin(partialProduct_5[7]));
wire wire_82, wire_83;
bit_adder add38(.S(wire_82), .Cout(wire_83),  .A(partialProduct_3[10]), .B(partialProduct_4[9]), .Cin(partialProduct_5[8]));
wire wire_84, wire_85;
bit_adder add39(.S(wire_84), .Cout(wire_85),  .A(partialProduct_3[11]), .B(partialProduct_4[10]), .Cin(partialProduct_5[9]));
wire wire_86, wire_87;
bit_adder add40(.S(wire_86), .Cout(wire_87),  .A(partialProduct_3[12]), .B(partialProduct_4[11]), .Cin(partialProduct_5[10]));
wire wire_88, wire_89;
bit_adder add41(.S(wire_88), .Cout(wire_89),  .A(partialProduct_3[13]), .B(partialProduct_4[12]), .Cin(partialProduct_5[11]));
wire wire_90, wire_91;
bit_adder add42(.S(wire_90), .Cout(wire_91),  .A(partialProduct_3[14]), .B(partialProduct_4[13]), .Cin(partialProduct_5[12]));
wire wire_92, wire_93;
bit_adder add43(.S(wire_92), .Cout(wire_93),  .A(partialProduct_3[15]), .B(partialProduct_4[14]), .Cin(partialProduct_5[13]));
wire wire_94, wire_95;
bit_adder add44(.S(wire_94), .Cout(wire_95),  .A(partialProduct_3[16]), .B(partialProduct_4[15]), .Cin(partialProduct_5[14]));
wire wire_96, wire_97;
bit_adder add45(.S(wire_96), .Cout(wire_97),  .A(partialProduct_3[17]), .B(partialProduct_4[16]), .Cin(partialProduct_5[15]));
wire wire_98, wire_99;
bit_adder add46(.S(wire_98), .Cout(wire_99),  .A(partialProduct_3[18]), .B(partialProduct_4[17]), .Cin(partialProduct_5[16]));
wire wire_100, wire_101;
bit_adder add47(.S(wire_100), .Cout(wire_101),  .A(partialProduct_3[19]), .B(partialProduct_4[18]), .Cin(partialProduct_5[17]));
wire wire_102, wire_103;
bit_adder add48(.S(wire_102), .Cout(wire_103),  .A(partialProduct_3[20]), .B(partialProduct_4[19]), .Cin(partialProduct_5[18]));
wire wire_104, wire_105;
bit_adder add49(.S(wire_104), .Cout(wire_105),  .A(partialProduct_3[21]), .B(partialProduct_4[20]), .Cin(partialProduct_5[19]));
wire wire_106, wire_107;
bit_adder add50(.S(wire_106), .Cout(wire_107),  .A(partialProduct_3[22]), .B(partialProduct_4[21]), .Cin(partialProduct_5[20]));
wire wire_108, wire_109;
bit_adder add51(.S(wire_108), .Cout(wire_109),  .A(partialProduct_3[23]), .B(partialProduct_4[22]), .Cin(partialProduct_5[21]));
wire wire_110, wire_111;
bit_adder add52(.S(wire_110), .Cout(wire_111),  .A(partialProduct_3[24]), .B(partialProduct_4[23]), .Cin(partialProduct_5[22]));
wire wire_112, wire_113;
bit_adder add53(.S(wire_112), .Cout(wire_113),  .A(partialProduct_3[25]), .B(partialProduct_4[24]), .Cin(partialProduct_5[23]));
wire wire_114, wire_115;
bit_adder add54(.S(wire_114), .Cout(wire_115),  .A(partialProduct_3[26]), .B(partialProduct_4[25]), .Cin(partialProduct_5[24]));
wire wire_116, wire_117;
bit_adder add55(.S(wire_116), .Cout(wire_117),  .A(partialProduct_3[27]), .B(partialProduct_4[26]), .Cin(partialProduct_5[25]));
wire wire_118, wire_119;
bit_adder add56(.S(wire_118), .Cout(wire_119),  .A(partialProduct_3[28]), .B(partialProduct_4[27]), .Cin(partialProduct_5[26]));
wire wire_120, wire_121;
bit_adder add57(.S(wire_120), .Cout(wire_121),  .A(partialProduct_3[29]), .B(partialProduct_4[28]), .Cin(partialProduct_5[27]));
wire wire_122, wire_123;
bit_adder add58(.S(wire_122), .Cout(wire_123),  .A(partialProduct_3[30]), .B(partialProduct_4[29]), .Cin(partialProduct_5[28]));
wire wire_124, wire_125;
bit_adder add59(.S(wire_124), .Cout(wire_125),  .A(partialProduct_3[31]), .B(partialProduct_4[30]), .Cin(partialProduct_5[29]));
wire wire_126, wire_127;
assign wire_126 = partialProduct_4[31] ^ partialProduct_5[30];
assign wire_127 = partialProduct_4[31] & partialProduct_5[30];
wire wire_128, wire_129;
assign wire_128 = partialProduct_6[1] ^ partialProduct_7[0];
assign wire_129 = partialProduct_6[1] & partialProduct_7[0];
wire wire_130, wire_131;
bit_adder add60(.S(wire_130), .Cout(wire_131),  .A(partialProduct_6[2]), .B(partialProduct_7[1]), .Cin(partialProduct_8[0]));
wire wire_132, wire_133;
bit_adder add61(.S(wire_132), .Cout(wire_133),  .A(partialProduct_6[3]), .B(partialProduct_7[2]), .Cin(partialProduct_8[1]));
wire wire_134, wire_135;
bit_adder add62(.S(wire_134), .Cout(wire_135),  .A(partialProduct_6[4]), .B(partialProduct_7[3]), .Cin(partialProduct_8[2]));
wire wire_136, wire_137;
bit_adder add63(.S(wire_136), .Cout(wire_137),  .A(partialProduct_6[5]), .B(partialProduct_7[4]), .Cin(partialProduct_8[3]));
wire wire_138, wire_139;
bit_adder add64(.S(wire_138), .Cout(wire_139),  .A(partialProduct_6[6]), .B(partialProduct_7[5]), .Cin(partialProduct_8[4]));
wire wire_140, wire_141;
bit_adder add65(.S(wire_140), .Cout(wire_141),  .A(partialProduct_6[7]), .B(partialProduct_7[6]), .Cin(partialProduct_8[5]));
wire wire_142, wire_143;
bit_adder add66(.S(wire_142), .Cout(wire_143),  .A(partialProduct_6[8]), .B(partialProduct_7[7]), .Cin(partialProduct_8[6]));
wire wire_144, wire_145;
bit_adder add67(.S(wire_144), .Cout(wire_145),  .A(partialProduct_6[9]), .B(partialProduct_7[8]), .Cin(partialProduct_8[7]));
wire wire_146, wire_147;
bit_adder add68(.S(wire_146), .Cout(wire_147),  .A(partialProduct_6[10]), .B(partialProduct_7[9]), .Cin(partialProduct_8[8]));
wire wire_148, wire_149;
bit_adder add69(.S(wire_148), .Cout(wire_149),  .A(partialProduct_6[11]), .B(partialProduct_7[10]), .Cin(partialProduct_8[9]));
wire wire_150, wire_151;
bit_adder add70(.S(wire_150), .Cout(wire_151),  .A(partialProduct_6[12]), .B(partialProduct_7[11]), .Cin(partialProduct_8[10]));
wire wire_152, wire_153;
bit_adder add71(.S(wire_152), .Cout(wire_153),  .A(partialProduct_6[13]), .B(partialProduct_7[12]), .Cin(partialProduct_8[11]));
wire wire_154, wire_155;
bit_adder add72(.S(wire_154), .Cout(wire_155),  .A(partialProduct_6[14]), .B(partialProduct_7[13]), .Cin(partialProduct_8[12]));
wire wire_156, wire_157;
bit_adder add73(.S(wire_156), .Cout(wire_157),  .A(partialProduct_6[15]), .B(partialProduct_7[14]), .Cin(partialProduct_8[13]));
wire wire_158, wire_159;
bit_adder add74(.S(wire_158), .Cout(wire_159),  .A(partialProduct_6[16]), .B(partialProduct_7[15]), .Cin(partialProduct_8[14]));
wire wire_160, wire_161;
bit_adder add75(.S(wire_160), .Cout(wire_161),  .A(partialProduct_6[17]), .B(partialProduct_7[16]), .Cin(partialProduct_8[15]));
wire wire_162, wire_163;
bit_adder add76(.S(wire_162), .Cout(wire_163),  .A(partialProduct_6[18]), .B(partialProduct_7[17]), .Cin(partialProduct_8[16]));
wire wire_164, wire_165;
bit_adder add77(.S(wire_164), .Cout(wire_165),  .A(partialProduct_6[19]), .B(partialProduct_7[18]), .Cin(partialProduct_8[17]));
wire wire_166, wire_167;
bit_adder add78(.S(wire_166), .Cout(wire_167),  .A(partialProduct_6[20]), .B(partialProduct_7[19]), .Cin(partialProduct_8[18]));
wire wire_168, wire_169;
bit_adder add79(.S(wire_168), .Cout(wire_169),  .A(partialProduct_6[21]), .B(partialProduct_7[20]), .Cin(partialProduct_8[19]));
wire wire_170, wire_171;
bit_adder add80(.S(wire_170), .Cout(wire_171),  .A(partialProduct_6[22]), .B(partialProduct_7[21]), .Cin(partialProduct_8[20]));
wire wire_172, wire_173;
bit_adder add81(.S(wire_172), .Cout(wire_173),  .A(partialProduct_6[23]), .B(partialProduct_7[22]), .Cin(partialProduct_8[21]));
wire wire_174, wire_175;
bit_adder add82(.S(wire_174), .Cout(wire_175),  .A(partialProduct_6[24]), .B(partialProduct_7[23]), .Cin(partialProduct_8[22]));
wire wire_176, wire_177;
bit_adder add83(.S(wire_176), .Cout(wire_177),  .A(partialProduct_6[25]), .B(partialProduct_7[24]), .Cin(partialProduct_8[23]));
wire wire_178, wire_179;
bit_adder add84(.S(wire_178), .Cout(wire_179),  .A(partialProduct_6[26]), .B(partialProduct_7[25]), .Cin(partialProduct_8[24]));
wire wire_180, wire_181;
bit_adder add85(.S(wire_180), .Cout(wire_181),  .A(partialProduct_6[27]), .B(partialProduct_7[26]), .Cin(partialProduct_8[25]));
wire wire_182, wire_183;
bit_adder add86(.S(wire_182), .Cout(wire_183),  .A(partialProduct_6[28]), .B(partialProduct_7[27]), .Cin(partialProduct_8[26]));
wire wire_184, wire_185;
bit_adder add87(.S(wire_184), .Cout(wire_185),  .A(partialProduct_6[29]), .B(partialProduct_7[28]), .Cin(partialProduct_8[27]));
wire wire_186, wire_187;
bit_adder add88(.S(wire_186), .Cout(wire_187),  .A(partialProduct_6[30]), .B(partialProduct_7[29]), .Cin(partialProduct_8[28]));
wire wire_188, wire_189;
bit_adder add89(.S(wire_188), .Cout(wire_189),  .A(partialProduct_6[31]), .B(partialProduct_7[30]), .Cin(partialProduct_8[29]));
wire wire_190, wire_191;
assign wire_190 = partialProduct_7[31] ^ partialProduct_8[30];
assign wire_191 = partialProduct_7[31] & partialProduct_8[30];
wire wire_192, wire_193;
assign wire_192 = partialProduct_9[1] ^ partialProduct_10[0];
assign wire_193 = partialProduct_9[1] & partialProduct_10[0];
wire wire_194, wire_195;
bit_adder add90(.S(wire_194), .Cout(wire_195),  .A(partialProduct_9[2]), .B(partialProduct_10[1]), .Cin(partialProduct_11[0]));
wire wire_196, wire_197;
bit_adder add91(.S(wire_196), .Cout(wire_197),  .A(partialProduct_9[3]), .B(partialProduct_10[2]), .Cin(partialProduct_11[1]));
wire wire_198, wire_199;
bit_adder add92(.S(wire_198), .Cout(wire_199),  .A(partialProduct_9[4]), .B(partialProduct_10[3]), .Cin(partialProduct_11[2]));
wire wire_200, wire_201;
bit_adder add93(.S(wire_200), .Cout(wire_201),  .A(partialProduct_9[5]), .B(partialProduct_10[4]), .Cin(partialProduct_11[3]));
wire wire_202, wire_203;
bit_adder add94(.S(wire_202), .Cout(wire_203),  .A(partialProduct_9[6]), .B(partialProduct_10[5]), .Cin(partialProduct_11[4]));
wire wire_204, wire_205;
bit_adder add95(.S(wire_204), .Cout(wire_205),  .A(partialProduct_9[7]), .B(partialProduct_10[6]), .Cin(partialProduct_11[5]));
wire wire_206, wire_207;
bit_adder add96(.S(wire_206), .Cout(wire_207),  .A(partialProduct_9[8]), .B(partialProduct_10[7]), .Cin(partialProduct_11[6]));
wire wire_208, wire_209;
bit_adder add97(.S(wire_208), .Cout(wire_209),  .A(partialProduct_9[9]), .B(partialProduct_10[8]), .Cin(partialProduct_11[7]));
wire wire_210, wire_211;
bit_adder add98(.S(wire_210), .Cout(wire_211),  .A(partialProduct_9[10]), .B(partialProduct_10[9]), .Cin(partialProduct_11[8]));
wire wire_212, wire_213;
bit_adder add99(.S(wire_212), .Cout(wire_213),  .A(partialProduct_9[11]), .B(partialProduct_10[10]), .Cin(partialProduct_11[9]));
wire wire_214, wire_215;
bit_adder add100(.S(wire_214), .Cout(wire_215),  .A(partialProduct_9[12]), .B(partialProduct_10[11]), .Cin(partialProduct_11[10]));
wire wire_216, wire_217;
bit_adder add101(.S(wire_216), .Cout(wire_217),  .A(partialProduct_9[13]), .B(partialProduct_10[12]), .Cin(partialProduct_11[11]));
wire wire_218, wire_219;
bit_adder add102(.S(wire_218), .Cout(wire_219),  .A(partialProduct_9[14]), .B(partialProduct_10[13]), .Cin(partialProduct_11[12]));
wire wire_220, wire_221;
bit_adder add103(.S(wire_220), .Cout(wire_221),  .A(partialProduct_9[15]), .B(partialProduct_10[14]), .Cin(partialProduct_11[13]));
wire wire_222, wire_223;
bit_adder add104(.S(wire_222), .Cout(wire_223),  .A(partialProduct_9[16]), .B(partialProduct_10[15]), .Cin(partialProduct_11[14]));
wire wire_224, wire_225;
bit_adder add105(.S(wire_224), .Cout(wire_225),  .A(partialProduct_9[17]), .B(partialProduct_10[16]), .Cin(partialProduct_11[15]));
wire wire_226, wire_227;
bit_adder add106(.S(wire_226), .Cout(wire_227),  .A(partialProduct_9[18]), .B(partialProduct_10[17]), .Cin(partialProduct_11[16]));
wire wire_228, wire_229;
bit_adder add107(.S(wire_228), .Cout(wire_229),  .A(partialProduct_9[19]), .B(partialProduct_10[18]), .Cin(partialProduct_11[17]));
wire wire_230, wire_231;
bit_adder add108(.S(wire_230), .Cout(wire_231),  .A(partialProduct_9[20]), .B(partialProduct_10[19]), .Cin(partialProduct_11[18]));
wire wire_232, wire_233;
bit_adder add109(.S(wire_232), .Cout(wire_233),  .A(partialProduct_9[21]), .B(partialProduct_10[20]), .Cin(partialProduct_11[19]));
wire wire_234, wire_235;
bit_adder add110(.S(wire_234), .Cout(wire_235),  .A(partialProduct_9[22]), .B(partialProduct_10[21]), .Cin(partialProduct_11[20]));
wire wire_236, wire_237;
bit_adder add111(.S(wire_236), .Cout(wire_237),  .A(partialProduct_9[23]), .B(partialProduct_10[22]), .Cin(partialProduct_11[21]));
wire wire_238, wire_239;
bit_adder add112(.S(wire_238), .Cout(wire_239),  .A(partialProduct_9[24]), .B(partialProduct_10[23]), .Cin(partialProduct_11[22]));
wire wire_240, wire_241;
bit_adder add113(.S(wire_240), .Cout(wire_241),  .A(partialProduct_9[25]), .B(partialProduct_10[24]), .Cin(partialProduct_11[23]));
wire wire_242, wire_243;
bit_adder add114(.S(wire_242), .Cout(wire_243),  .A(partialProduct_9[26]), .B(partialProduct_10[25]), .Cin(partialProduct_11[24]));
wire wire_244, wire_245;
bit_adder add115(.S(wire_244), .Cout(wire_245),  .A(partialProduct_9[27]), .B(partialProduct_10[26]), .Cin(partialProduct_11[25]));
wire wire_246, wire_247;
bit_adder add116(.S(wire_246), .Cout(wire_247),  .A(partialProduct_9[28]), .B(partialProduct_10[27]), .Cin(partialProduct_11[26]));
wire wire_248, wire_249;
bit_adder add117(.S(wire_248), .Cout(wire_249),  .A(partialProduct_9[29]), .B(partialProduct_10[28]), .Cin(partialProduct_11[27]));
wire wire_250, wire_251;
bit_adder add118(.S(wire_250), .Cout(wire_251),  .A(partialProduct_9[30]), .B(partialProduct_10[29]), .Cin(partialProduct_11[28]));
wire wire_252, wire_253;
bit_adder add119(.S(wire_252), .Cout(wire_253),  .A(partialProduct_9[31]), .B(partialProduct_10[30]), .Cin(partialProduct_11[29]));
wire wire_254, wire_255;
assign wire_254 = partialProduct_10[31] ^ partialProduct_11[30];
assign wire_255 = partialProduct_10[31] & partialProduct_11[30];
wire wire_256, wire_257;
assign wire_256 = partialProduct_12[1] ^ partialProduct_13[0];
assign wire_257 = partialProduct_12[1] & partialProduct_13[0];
wire wire_258, wire_259;
bit_adder add120(.S(wire_258), .Cout(wire_259),  .A(partialProduct_12[2]), .B(partialProduct_13[1]), .Cin(partialProduct_14[0]));
wire wire_260, wire_261;
bit_adder add121(.S(wire_260), .Cout(wire_261),  .A(partialProduct_12[3]), .B(partialProduct_13[2]), .Cin(partialProduct_14[1]));
wire wire_262, wire_263;
bit_adder add122(.S(wire_262), .Cout(wire_263),  .A(partialProduct_12[4]), .B(partialProduct_13[3]), .Cin(partialProduct_14[2]));
wire wire_264, wire_265;
bit_adder add123(.S(wire_264), .Cout(wire_265),  .A(partialProduct_12[5]), .B(partialProduct_13[4]), .Cin(partialProduct_14[3]));
wire wire_266, wire_267;
bit_adder add124(.S(wire_266), .Cout(wire_267),  .A(partialProduct_12[6]), .B(partialProduct_13[5]), .Cin(partialProduct_14[4]));
wire wire_268, wire_269;
bit_adder add125(.S(wire_268), .Cout(wire_269),  .A(partialProduct_12[7]), .B(partialProduct_13[6]), .Cin(partialProduct_14[5]));
wire wire_270, wire_271;
bit_adder add126(.S(wire_270), .Cout(wire_271),  .A(partialProduct_12[8]), .B(partialProduct_13[7]), .Cin(partialProduct_14[6]));
wire wire_272, wire_273;
bit_adder add127(.S(wire_272), .Cout(wire_273),  .A(partialProduct_12[9]), .B(partialProduct_13[8]), .Cin(partialProduct_14[7]));
wire wire_274, wire_275;
bit_adder add128(.S(wire_274), .Cout(wire_275),  .A(partialProduct_12[10]), .B(partialProduct_13[9]), .Cin(partialProduct_14[8]));
wire wire_276, wire_277;
bit_adder add129(.S(wire_276), .Cout(wire_277),  .A(partialProduct_12[11]), .B(partialProduct_13[10]), .Cin(partialProduct_14[9]));
wire wire_278, wire_279;
bit_adder add130(.S(wire_278), .Cout(wire_279),  .A(partialProduct_12[12]), .B(partialProduct_13[11]), .Cin(partialProduct_14[10]));
wire wire_280, wire_281;
bit_adder add131(.S(wire_280), .Cout(wire_281),  .A(partialProduct_12[13]), .B(partialProduct_13[12]), .Cin(partialProduct_14[11]));
wire wire_282, wire_283;
bit_adder add132(.S(wire_282), .Cout(wire_283),  .A(partialProduct_12[14]), .B(partialProduct_13[13]), .Cin(partialProduct_14[12]));
wire wire_284, wire_285;
bit_adder add133(.S(wire_284), .Cout(wire_285),  .A(partialProduct_12[15]), .B(partialProduct_13[14]), .Cin(partialProduct_14[13]));
wire wire_286, wire_287;
bit_adder add134(.S(wire_286), .Cout(wire_287),  .A(partialProduct_12[16]), .B(partialProduct_13[15]), .Cin(partialProduct_14[14]));
wire wire_288, wire_289;
bit_adder add135(.S(wire_288), .Cout(wire_289),  .A(partialProduct_12[17]), .B(partialProduct_13[16]), .Cin(partialProduct_14[15]));
wire wire_290, wire_291;
bit_adder add136(.S(wire_290), .Cout(wire_291),  .A(partialProduct_12[18]), .B(partialProduct_13[17]), .Cin(partialProduct_14[16]));
wire wire_292, wire_293;
bit_adder add137(.S(wire_292), .Cout(wire_293),  .A(partialProduct_12[19]), .B(partialProduct_13[18]), .Cin(partialProduct_14[17]));
wire wire_294, wire_295;
bit_adder add138(.S(wire_294), .Cout(wire_295),  .A(partialProduct_12[20]), .B(partialProduct_13[19]), .Cin(partialProduct_14[18]));
wire wire_296, wire_297;
bit_adder add139(.S(wire_296), .Cout(wire_297),  .A(partialProduct_12[21]), .B(partialProduct_13[20]), .Cin(partialProduct_14[19]));
wire wire_298, wire_299;
bit_adder add140(.S(wire_298), .Cout(wire_299),  .A(partialProduct_12[22]), .B(partialProduct_13[21]), .Cin(partialProduct_14[20]));
wire wire_300, wire_301;
bit_adder add141(.S(wire_300), .Cout(wire_301),  .A(partialProduct_12[23]), .B(partialProduct_13[22]), .Cin(partialProduct_14[21]));
wire wire_302, wire_303;
bit_adder add142(.S(wire_302), .Cout(wire_303),  .A(partialProduct_12[24]), .B(partialProduct_13[23]), .Cin(partialProduct_14[22]));
wire wire_304, wire_305;
bit_adder add143(.S(wire_304), .Cout(wire_305),  .A(partialProduct_12[25]), .B(partialProduct_13[24]), .Cin(partialProduct_14[23]));
wire wire_306, wire_307;
bit_adder add144(.S(wire_306), .Cout(wire_307),  .A(partialProduct_12[26]), .B(partialProduct_13[25]), .Cin(partialProduct_14[24]));
wire wire_308, wire_309;
bit_adder add145(.S(wire_308), .Cout(wire_309),  .A(partialProduct_12[27]), .B(partialProduct_13[26]), .Cin(partialProduct_14[25]));
wire wire_310, wire_311;
bit_adder add146(.S(wire_310), .Cout(wire_311),  .A(partialProduct_12[28]), .B(partialProduct_13[27]), .Cin(partialProduct_14[26]));
wire wire_312, wire_313;
bit_adder add147(.S(wire_312), .Cout(wire_313),  .A(partialProduct_12[29]), .B(partialProduct_13[28]), .Cin(partialProduct_14[27]));
wire wire_314, wire_315;
bit_adder add148(.S(wire_314), .Cout(wire_315),  .A(partialProduct_12[30]), .B(partialProduct_13[29]), .Cin(partialProduct_14[28]));
wire wire_316, wire_317;
bit_adder add149(.S(wire_316), .Cout(wire_317),  .A(partialProduct_12[31]), .B(partialProduct_13[30]), .Cin(partialProduct_14[29]));
wire wire_318, wire_319;
assign wire_318 = partialProduct_13[31] ^ partialProduct_14[30];
assign wire_319 = partialProduct_13[31] & partialProduct_14[30];
wire wire_320, wire_321;
assign wire_320 = partialProduct_15[1] ^ partialProduct_16[0];
assign wire_321 = partialProduct_15[1] & partialProduct_16[0];
wire wire_322, wire_323;
bit_adder add150(.S(wire_322), .Cout(wire_323),  .A(partialProduct_15[2]), .B(partialProduct_16[1]), .Cin(partialProduct_17[0]));
wire wire_324, wire_325;
bit_adder add151(.S(wire_324), .Cout(wire_325),  .A(partialProduct_15[3]), .B(partialProduct_16[2]), .Cin(partialProduct_17[1]));
wire wire_326, wire_327;
bit_adder add152(.S(wire_326), .Cout(wire_327),  .A(partialProduct_15[4]), .B(partialProduct_16[3]), .Cin(partialProduct_17[2]));
wire wire_328, wire_329;
bit_adder add153(.S(wire_328), .Cout(wire_329),  .A(partialProduct_15[5]), .B(partialProduct_16[4]), .Cin(partialProduct_17[3]));
wire wire_330, wire_331;
bit_adder add154(.S(wire_330), .Cout(wire_331),  .A(partialProduct_15[6]), .B(partialProduct_16[5]), .Cin(partialProduct_17[4]));
wire wire_332, wire_333;
bit_adder add155(.S(wire_332), .Cout(wire_333),  .A(partialProduct_15[7]), .B(partialProduct_16[6]), .Cin(partialProduct_17[5]));
wire wire_334, wire_335;
bit_adder add156(.S(wire_334), .Cout(wire_335),  .A(partialProduct_15[8]), .B(partialProduct_16[7]), .Cin(partialProduct_17[6]));
wire wire_336, wire_337;
bit_adder add157(.S(wire_336), .Cout(wire_337),  .A(partialProduct_15[9]), .B(partialProduct_16[8]), .Cin(partialProduct_17[7]));
wire wire_338, wire_339;
bit_adder add158(.S(wire_338), .Cout(wire_339),  .A(partialProduct_15[10]), .B(partialProduct_16[9]), .Cin(partialProduct_17[8]));
wire wire_340, wire_341;
bit_adder add159(.S(wire_340), .Cout(wire_341),  .A(partialProduct_15[11]), .B(partialProduct_16[10]), .Cin(partialProduct_17[9]));
wire wire_342, wire_343;
bit_adder add160(.S(wire_342), .Cout(wire_343),  .A(partialProduct_15[12]), .B(partialProduct_16[11]), .Cin(partialProduct_17[10]));
wire wire_344, wire_345;
bit_adder add161(.S(wire_344), .Cout(wire_345),  .A(partialProduct_15[13]), .B(partialProduct_16[12]), .Cin(partialProduct_17[11]));
wire wire_346, wire_347;
bit_adder add162(.S(wire_346), .Cout(wire_347),  .A(partialProduct_15[14]), .B(partialProduct_16[13]), .Cin(partialProduct_17[12]));
wire wire_348, wire_349;
bit_adder add163(.S(wire_348), .Cout(wire_349),  .A(partialProduct_15[15]), .B(partialProduct_16[14]), .Cin(partialProduct_17[13]));
wire wire_350, wire_351;
bit_adder add164(.S(wire_350), .Cout(wire_351),  .A(partialProduct_15[16]), .B(partialProduct_16[15]), .Cin(partialProduct_17[14]));
wire wire_352, wire_353;
bit_adder add165(.S(wire_352), .Cout(wire_353),  .A(partialProduct_15[17]), .B(partialProduct_16[16]), .Cin(partialProduct_17[15]));
wire wire_354, wire_355;
bit_adder add166(.S(wire_354), .Cout(wire_355),  .A(partialProduct_15[18]), .B(partialProduct_16[17]), .Cin(partialProduct_17[16]));
wire wire_356, wire_357;
bit_adder add167(.S(wire_356), .Cout(wire_357),  .A(partialProduct_15[19]), .B(partialProduct_16[18]), .Cin(partialProduct_17[17]));
wire wire_358, wire_359;
bit_adder add168(.S(wire_358), .Cout(wire_359),  .A(partialProduct_15[20]), .B(partialProduct_16[19]), .Cin(partialProduct_17[18]));
wire wire_360, wire_361;
bit_adder add169(.S(wire_360), .Cout(wire_361),  .A(partialProduct_15[21]), .B(partialProduct_16[20]), .Cin(partialProduct_17[19]));
wire wire_362, wire_363;
bit_adder add170(.S(wire_362), .Cout(wire_363),  .A(partialProduct_15[22]), .B(partialProduct_16[21]), .Cin(partialProduct_17[20]));
wire wire_364, wire_365;
bit_adder add171(.S(wire_364), .Cout(wire_365),  .A(partialProduct_15[23]), .B(partialProduct_16[22]), .Cin(partialProduct_17[21]));
wire wire_366, wire_367;
bit_adder add172(.S(wire_366), .Cout(wire_367),  .A(partialProduct_15[24]), .B(partialProduct_16[23]), .Cin(partialProduct_17[22]));
wire wire_368, wire_369;
bit_adder add173(.S(wire_368), .Cout(wire_369),  .A(partialProduct_15[25]), .B(partialProduct_16[24]), .Cin(partialProduct_17[23]));
wire wire_370, wire_371;
bit_adder add174(.S(wire_370), .Cout(wire_371),  .A(partialProduct_15[26]), .B(partialProduct_16[25]), .Cin(partialProduct_17[24]));
wire wire_372, wire_373;
bit_adder add175(.S(wire_372), .Cout(wire_373),  .A(partialProduct_15[27]), .B(partialProduct_16[26]), .Cin(partialProduct_17[25]));
wire wire_374, wire_375;
bit_adder add176(.S(wire_374), .Cout(wire_375),  .A(partialProduct_15[28]), .B(partialProduct_16[27]), .Cin(partialProduct_17[26]));
wire wire_376, wire_377;
bit_adder add177(.S(wire_376), .Cout(wire_377),  .A(partialProduct_15[29]), .B(partialProduct_16[28]), .Cin(partialProduct_17[27]));
wire wire_378, wire_379;
bit_adder add178(.S(wire_378), .Cout(wire_379),  .A(partialProduct_15[30]), .B(partialProduct_16[29]), .Cin(partialProduct_17[28]));
wire wire_380, wire_381;
bit_adder add179(.S(wire_380), .Cout(wire_381),  .A(partialProduct_15[31]), .B(partialProduct_16[30]), .Cin(partialProduct_17[29]));
wire wire_382, wire_383;
assign wire_382 = partialProduct_16[31] ^ partialProduct_17[30];
assign wire_383 = partialProduct_16[31] & partialProduct_17[30];
wire wire_384, wire_385;
assign wire_384 = partialProduct_18[1] ^ partialProduct_19[0];
assign wire_385 = partialProduct_18[1] & partialProduct_19[0];
wire wire_386, wire_387;
bit_adder add180(.S(wire_386), .Cout(wire_387),  .A(partialProduct_18[2]), .B(partialProduct_19[1]), .Cin(partialProduct_20[0]));
wire wire_388, wire_389;
bit_adder add181(.S(wire_388), .Cout(wire_389),  .A(partialProduct_18[3]), .B(partialProduct_19[2]), .Cin(partialProduct_20[1]));
wire wire_390, wire_391;
bit_adder add182(.S(wire_390), .Cout(wire_391),  .A(partialProduct_18[4]), .B(partialProduct_19[3]), .Cin(partialProduct_20[2]));
wire wire_392, wire_393;
bit_adder add183(.S(wire_392), .Cout(wire_393),  .A(partialProduct_18[5]), .B(partialProduct_19[4]), .Cin(partialProduct_20[3]));
wire wire_394, wire_395;
bit_adder add184(.S(wire_394), .Cout(wire_395),  .A(partialProduct_18[6]), .B(partialProduct_19[5]), .Cin(partialProduct_20[4]));
wire wire_396, wire_397;
bit_adder add185(.S(wire_396), .Cout(wire_397),  .A(partialProduct_18[7]), .B(partialProduct_19[6]), .Cin(partialProduct_20[5]));
wire wire_398, wire_399;
bit_adder add186(.S(wire_398), .Cout(wire_399),  .A(partialProduct_18[8]), .B(partialProduct_19[7]), .Cin(partialProduct_20[6]));
wire wire_400, wire_401;
bit_adder add187(.S(wire_400), .Cout(wire_401),  .A(partialProduct_18[9]), .B(partialProduct_19[8]), .Cin(partialProduct_20[7]));
wire wire_402, wire_403;
bit_adder add188(.S(wire_402), .Cout(wire_403),  .A(partialProduct_18[10]), .B(partialProduct_19[9]), .Cin(partialProduct_20[8]));
wire wire_404, wire_405;
bit_adder add189(.S(wire_404), .Cout(wire_405),  .A(partialProduct_18[11]), .B(partialProduct_19[10]), .Cin(partialProduct_20[9]));
wire wire_406, wire_407;
bit_adder add190(.S(wire_406), .Cout(wire_407),  .A(partialProduct_18[12]), .B(partialProduct_19[11]), .Cin(partialProduct_20[10]));
wire wire_408, wire_409;
bit_adder add191(.S(wire_408), .Cout(wire_409),  .A(partialProduct_18[13]), .B(partialProduct_19[12]), .Cin(partialProduct_20[11]));
wire wire_410, wire_411;
bit_adder add192(.S(wire_410), .Cout(wire_411),  .A(partialProduct_18[14]), .B(partialProduct_19[13]), .Cin(partialProduct_20[12]));
wire wire_412, wire_413;
bit_adder add193(.S(wire_412), .Cout(wire_413),  .A(partialProduct_18[15]), .B(partialProduct_19[14]), .Cin(partialProduct_20[13]));
wire wire_414, wire_415;
bit_adder add194(.S(wire_414), .Cout(wire_415),  .A(partialProduct_18[16]), .B(partialProduct_19[15]), .Cin(partialProduct_20[14]));
wire wire_416, wire_417;
bit_adder add195(.S(wire_416), .Cout(wire_417),  .A(partialProduct_18[17]), .B(partialProduct_19[16]), .Cin(partialProduct_20[15]));
wire wire_418, wire_419;
bit_adder add196(.S(wire_418), .Cout(wire_419),  .A(partialProduct_18[18]), .B(partialProduct_19[17]), .Cin(partialProduct_20[16]));
wire wire_420, wire_421;
bit_adder add197(.S(wire_420), .Cout(wire_421),  .A(partialProduct_18[19]), .B(partialProduct_19[18]), .Cin(partialProduct_20[17]));
wire wire_422, wire_423;
bit_adder add198(.S(wire_422), .Cout(wire_423),  .A(partialProduct_18[20]), .B(partialProduct_19[19]), .Cin(partialProduct_20[18]));
wire wire_424, wire_425;
bit_adder add199(.S(wire_424), .Cout(wire_425),  .A(partialProduct_18[21]), .B(partialProduct_19[20]), .Cin(partialProduct_20[19]));
wire wire_426, wire_427;
bit_adder add200(.S(wire_426), .Cout(wire_427),  .A(partialProduct_18[22]), .B(partialProduct_19[21]), .Cin(partialProduct_20[20]));
wire wire_428, wire_429;
bit_adder add201(.S(wire_428), .Cout(wire_429),  .A(partialProduct_18[23]), .B(partialProduct_19[22]), .Cin(partialProduct_20[21]));
wire wire_430, wire_431;
bit_adder add202(.S(wire_430), .Cout(wire_431),  .A(partialProduct_18[24]), .B(partialProduct_19[23]), .Cin(partialProduct_20[22]));
wire wire_432, wire_433;
bit_adder add203(.S(wire_432), .Cout(wire_433),  .A(partialProduct_18[25]), .B(partialProduct_19[24]), .Cin(partialProduct_20[23]));
wire wire_434, wire_435;
bit_adder add204(.S(wire_434), .Cout(wire_435),  .A(partialProduct_18[26]), .B(partialProduct_19[25]), .Cin(partialProduct_20[24]));
wire wire_436, wire_437;
bit_adder add205(.S(wire_436), .Cout(wire_437),  .A(partialProduct_18[27]), .B(partialProduct_19[26]), .Cin(partialProduct_20[25]));
wire wire_438, wire_439;
bit_adder add206(.S(wire_438), .Cout(wire_439),  .A(partialProduct_18[28]), .B(partialProduct_19[27]), .Cin(partialProduct_20[26]));
wire wire_440, wire_441;
bit_adder add207(.S(wire_440), .Cout(wire_441),  .A(partialProduct_18[29]), .B(partialProduct_19[28]), .Cin(partialProduct_20[27]));
wire wire_442, wire_443;
bit_adder add208(.S(wire_442), .Cout(wire_443),  .A(partialProduct_18[30]), .B(partialProduct_19[29]), .Cin(partialProduct_20[28]));
wire wire_444, wire_445;
bit_adder add209(.S(wire_444), .Cout(wire_445),  .A(partialProduct_18[31]), .B(partialProduct_19[30]), .Cin(partialProduct_20[29]));
wire wire_446, wire_447;
assign wire_446 = partialProduct_19[31] ^ partialProduct_20[30];
assign wire_447 = partialProduct_19[31] & partialProduct_20[30];
wire wire_448, wire_449;
assign wire_448 = partialProduct_21[1] ^ partialProduct_22[0];
assign wire_449 = partialProduct_21[1] & partialProduct_22[0];
wire wire_450, wire_451;
bit_adder add210(.S(wire_450), .Cout(wire_451),  .A(partialProduct_21[2]), .B(partialProduct_22[1]), .Cin(partialProduct_23[0]));
wire wire_452, wire_453;
bit_adder add211(.S(wire_452), .Cout(wire_453),  .A(partialProduct_21[3]), .B(partialProduct_22[2]), .Cin(partialProduct_23[1]));
wire wire_454, wire_455;
bit_adder add212(.S(wire_454), .Cout(wire_455),  .A(partialProduct_21[4]), .B(partialProduct_22[3]), .Cin(partialProduct_23[2]));
wire wire_456, wire_457;
bit_adder add213(.S(wire_456), .Cout(wire_457),  .A(partialProduct_21[5]), .B(partialProduct_22[4]), .Cin(partialProduct_23[3]));
wire wire_458, wire_459;
bit_adder add214(.S(wire_458), .Cout(wire_459),  .A(partialProduct_21[6]), .B(partialProduct_22[5]), .Cin(partialProduct_23[4]));
wire wire_460, wire_461;
bit_adder add215(.S(wire_460), .Cout(wire_461),  .A(partialProduct_21[7]), .B(partialProduct_22[6]), .Cin(partialProduct_23[5]));
wire wire_462, wire_463;
bit_adder add216(.S(wire_462), .Cout(wire_463),  .A(partialProduct_21[8]), .B(partialProduct_22[7]), .Cin(partialProduct_23[6]));
wire wire_464, wire_465;
bit_adder add217(.S(wire_464), .Cout(wire_465),  .A(partialProduct_21[9]), .B(partialProduct_22[8]), .Cin(partialProduct_23[7]));
wire wire_466, wire_467;
bit_adder add218(.S(wire_466), .Cout(wire_467),  .A(partialProduct_21[10]), .B(partialProduct_22[9]), .Cin(partialProduct_23[8]));
wire wire_468, wire_469;
bit_adder add219(.S(wire_468), .Cout(wire_469),  .A(partialProduct_21[11]), .B(partialProduct_22[10]), .Cin(partialProduct_23[9]));
wire wire_470, wire_471;
bit_adder add220(.S(wire_470), .Cout(wire_471),  .A(partialProduct_21[12]), .B(partialProduct_22[11]), .Cin(partialProduct_23[10]));
wire wire_472, wire_473;
bit_adder add221(.S(wire_472), .Cout(wire_473),  .A(partialProduct_21[13]), .B(partialProduct_22[12]), .Cin(partialProduct_23[11]));
wire wire_474, wire_475;
bit_adder add222(.S(wire_474), .Cout(wire_475),  .A(partialProduct_21[14]), .B(partialProduct_22[13]), .Cin(partialProduct_23[12]));
wire wire_476, wire_477;
bit_adder add223(.S(wire_476), .Cout(wire_477),  .A(partialProduct_21[15]), .B(partialProduct_22[14]), .Cin(partialProduct_23[13]));
wire wire_478, wire_479;
bit_adder add224(.S(wire_478), .Cout(wire_479),  .A(partialProduct_21[16]), .B(partialProduct_22[15]), .Cin(partialProduct_23[14]));
wire wire_480, wire_481;
bit_adder add225(.S(wire_480), .Cout(wire_481),  .A(partialProduct_21[17]), .B(partialProduct_22[16]), .Cin(partialProduct_23[15]));
wire wire_482, wire_483;
bit_adder add226(.S(wire_482), .Cout(wire_483),  .A(partialProduct_21[18]), .B(partialProduct_22[17]), .Cin(partialProduct_23[16]));
wire wire_484, wire_485;
bit_adder add227(.S(wire_484), .Cout(wire_485),  .A(partialProduct_21[19]), .B(partialProduct_22[18]), .Cin(partialProduct_23[17]));
wire wire_486, wire_487;
bit_adder add228(.S(wire_486), .Cout(wire_487),  .A(partialProduct_21[20]), .B(partialProduct_22[19]), .Cin(partialProduct_23[18]));
wire wire_488, wire_489;
bit_adder add229(.S(wire_488), .Cout(wire_489),  .A(partialProduct_21[21]), .B(partialProduct_22[20]), .Cin(partialProduct_23[19]));
wire wire_490, wire_491;
bit_adder add230(.S(wire_490), .Cout(wire_491),  .A(partialProduct_21[22]), .B(partialProduct_22[21]), .Cin(partialProduct_23[20]));
wire wire_492, wire_493;
bit_adder add231(.S(wire_492), .Cout(wire_493),  .A(partialProduct_21[23]), .B(partialProduct_22[22]), .Cin(partialProduct_23[21]));
wire wire_494, wire_495;
bit_adder add232(.S(wire_494), .Cout(wire_495),  .A(partialProduct_21[24]), .B(partialProduct_22[23]), .Cin(partialProduct_23[22]));
wire wire_496, wire_497;
bit_adder add233(.S(wire_496), .Cout(wire_497),  .A(partialProduct_21[25]), .B(partialProduct_22[24]), .Cin(partialProduct_23[23]));
wire wire_498, wire_499;
bit_adder add234(.S(wire_498), .Cout(wire_499),  .A(partialProduct_21[26]), .B(partialProduct_22[25]), .Cin(partialProduct_23[24]));
wire wire_500, wire_501;
bit_adder add235(.S(wire_500), .Cout(wire_501),  .A(partialProduct_21[27]), .B(partialProduct_22[26]), .Cin(partialProduct_23[25]));
wire wire_502, wire_503;
bit_adder add236(.S(wire_502), .Cout(wire_503),  .A(partialProduct_21[28]), .B(partialProduct_22[27]), .Cin(partialProduct_23[26]));
wire wire_504, wire_505;
bit_adder add237(.S(wire_504), .Cout(wire_505),  .A(partialProduct_21[29]), .B(partialProduct_22[28]), .Cin(partialProduct_23[27]));
wire wire_506, wire_507;
bit_adder add238(.S(wire_506), .Cout(wire_507),  .A(partialProduct_21[30]), .B(partialProduct_22[29]), .Cin(partialProduct_23[28]));
wire wire_508, wire_509;
bit_adder add239(.S(wire_508), .Cout(wire_509),  .A(partialProduct_21[31]), .B(partialProduct_22[30]), .Cin(partialProduct_23[29]));
wire wire_510, wire_511;
assign wire_510 = partialProduct_22[31] ^ partialProduct_23[30];
assign wire_511 = partialProduct_22[31] & partialProduct_23[30];
wire wire_512, wire_513;
assign wire_512 = partialProduct_24[1] ^ partialProduct_25[0];
assign wire_513 = partialProduct_24[1] & partialProduct_25[0];
wire wire_514, wire_515;
bit_adder add240(.S(wire_514), .Cout(wire_515),  .A(partialProduct_24[2]), .B(partialProduct_25[1]), .Cin(partialProduct_26[0]));
wire wire_516, wire_517;
bit_adder add241(.S(wire_516), .Cout(wire_517),  .A(partialProduct_24[3]), .B(partialProduct_25[2]), .Cin(partialProduct_26[1]));
wire wire_518, wire_519;
bit_adder add242(.S(wire_518), .Cout(wire_519),  .A(partialProduct_24[4]), .B(partialProduct_25[3]), .Cin(partialProduct_26[2]));
wire wire_520, wire_521;
bit_adder add243(.S(wire_520), .Cout(wire_521),  .A(partialProduct_24[5]), .B(partialProduct_25[4]), .Cin(partialProduct_26[3]));
wire wire_522, wire_523;
bit_adder add244(.S(wire_522), .Cout(wire_523),  .A(partialProduct_24[6]), .B(partialProduct_25[5]), .Cin(partialProduct_26[4]));
wire wire_524, wire_525;
bit_adder add245(.S(wire_524), .Cout(wire_525),  .A(partialProduct_24[7]), .B(partialProduct_25[6]), .Cin(partialProduct_26[5]));
wire wire_526, wire_527;
bit_adder add246(.S(wire_526), .Cout(wire_527),  .A(partialProduct_24[8]), .B(partialProduct_25[7]), .Cin(partialProduct_26[6]));
wire wire_528, wire_529;
bit_adder add247(.S(wire_528), .Cout(wire_529),  .A(partialProduct_24[9]), .B(partialProduct_25[8]), .Cin(partialProduct_26[7]));
wire wire_530, wire_531;
bit_adder add248(.S(wire_530), .Cout(wire_531),  .A(partialProduct_24[10]), .B(partialProduct_25[9]), .Cin(partialProduct_26[8]));
wire wire_532, wire_533;
bit_adder add249(.S(wire_532), .Cout(wire_533),  .A(partialProduct_24[11]), .B(partialProduct_25[10]), .Cin(partialProduct_26[9]));
wire wire_534, wire_535;
bit_adder add250(.S(wire_534), .Cout(wire_535),  .A(partialProduct_24[12]), .B(partialProduct_25[11]), .Cin(partialProduct_26[10]));
wire wire_536, wire_537;
bit_adder add251(.S(wire_536), .Cout(wire_537),  .A(partialProduct_24[13]), .B(partialProduct_25[12]), .Cin(partialProduct_26[11]));
wire wire_538, wire_539;
bit_adder add252(.S(wire_538), .Cout(wire_539),  .A(partialProduct_24[14]), .B(partialProduct_25[13]), .Cin(partialProduct_26[12]));
wire wire_540, wire_541;
bit_adder add253(.S(wire_540), .Cout(wire_541),  .A(partialProduct_24[15]), .B(partialProduct_25[14]), .Cin(partialProduct_26[13]));
wire wire_542, wire_543;
bit_adder add254(.S(wire_542), .Cout(wire_543),  .A(partialProduct_24[16]), .B(partialProduct_25[15]), .Cin(partialProduct_26[14]));
wire wire_544, wire_545;
bit_adder add255(.S(wire_544), .Cout(wire_545),  .A(partialProduct_24[17]), .B(partialProduct_25[16]), .Cin(partialProduct_26[15]));
wire wire_546, wire_547;
bit_adder add256(.S(wire_546), .Cout(wire_547),  .A(partialProduct_24[18]), .B(partialProduct_25[17]), .Cin(partialProduct_26[16]));
wire wire_548, wire_549;
bit_adder add257(.S(wire_548), .Cout(wire_549),  .A(partialProduct_24[19]), .B(partialProduct_25[18]), .Cin(partialProduct_26[17]));
wire wire_550, wire_551;
bit_adder add258(.S(wire_550), .Cout(wire_551),  .A(partialProduct_24[20]), .B(partialProduct_25[19]), .Cin(partialProduct_26[18]));
wire wire_552, wire_553;
bit_adder add259(.S(wire_552), .Cout(wire_553),  .A(partialProduct_24[21]), .B(partialProduct_25[20]), .Cin(partialProduct_26[19]));
wire wire_554, wire_555;
bit_adder add260(.S(wire_554), .Cout(wire_555),  .A(partialProduct_24[22]), .B(partialProduct_25[21]), .Cin(partialProduct_26[20]));
wire wire_556, wire_557;
bit_adder add261(.S(wire_556), .Cout(wire_557),  .A(partialProduct_24[23]), .B(partialProduct_25[22]), .Cin(partialProduct_26[21]));
wire wire_558, wire_559;
bit_adder add262(.S(wire_558), .Cout(wire_559),  .A(partialProduct_24[24]), .B(partialProduct_25[23]), .Cin(partialProduct_26[22]));
wire wire_560, wire_561;
bit_adder add263(.S(wire_560), .Cout(wire_561),  .A(partialProduct_24[25]), .B(partialProduct_25[24]), .Cin(partialProduct_26[23]));
wire wire_562, wire_563;
bit_adder add264(.S(wire_562), .Cout(wire_563),  .A(partialProduct_24[26]), .B(partialProduct_25[25]), .Cin(partialProduct_26[24]));
wire wire_564, wire_565;
bit_adder add265(.S(wire_564), .Cout(wire_565),  .A(partialProduct_24[27]), .B(partialProduct_25[26]), .Cin(partialProduct_26[25]));
wire wire_566, wire_567;
bit_adder add266(.S(wire_566), .Cout(wire_567),  .A(partialProduct_24[28]), .B(partialProduct_25[27]), .Cin(partialProduct_26[26]));
wire wire_568, wire_569;
bit_adder add267(.S(wire_568), .Cout(wire_569),  .A(partialProduct_24[29]), .B(partialProduct_25[28]), .Cin(partialProduct_26[27]));
wire wire_570, wire_571;
bit_adder add268(.S(wire_570), .Cout(wire_571),  .A(partialProduct_24[30]), .B(partialProduct_25[29]), .Cin(partialProduct_26[28]));
wire wire_572, wire_573;
bit_adder add269(.S(wire_572), .Cout(wire_573),  .A(partialProduct_24[31]), .B(partialProduct_25[30]), .Cin(partialProduct_26[29]));
wire wire_574, wire_575;
assign wire_574 = partialProduct_25[31] ^ partialProduct_26[30];
assign wire_575 = partialProduct_25[31] & partialProduct_26[30];
wire wire_576, wire_577;
assign wire_576 = partialProduct_27[1] ^ partialProduct_28[0];
assign wire_577 = partialProduct_27[1] & partialProduct_28[0];
wire wire_578, wire_579;
bit_adder add270(.S(wire_578), .Cout(wire_579),  .A(partialProduct_27[2]), .B(partialProduct_28[1]), .Cin(partialProduct_29[0]));
wire wire_580, wire_581;
bit_adder add271(.S(wire_580), .Cout(wire_581),  .A(partialProduct_27[3]), .B(partialProduct_28[2]), .Cin(partialProduct_29[1]));
wire wire_582, wire_583;
bit_adder add272(.S(wire_582), .Cout(wire_583),  .A(partialProduct_27[4]), .B(partialProduct_28[3]), .Cin(partialProduct_29[2]));
wire wire_584, wire_585;
bit_adder add273(.S(wire_584), .Cout(wire_585),  .A(partialProduct_27[5]), .B(partialProduct_28[4]), .Cin(partialProduct_29[3]));
wire wire_586, wire_587;
bit_adder add274(.S(wire_586), .Cout(wire_587),  .A(partialProduct_27[6]), .B(partialProduct_28[5]), .Cin(partialProduct_29[4]));
wire wire_588, wire_589;
bit_adder add275(.S(wire_588), .Cout(wire_589),  .A(partialProduct_27[7]), .B(partialProduct_28[6]), .Cin(partialProduct_29[5]));
wire wire_590, wire_591;
bit_adder add276(.S(wire_590), .Cout(wire_591),  .A(partialProduct_27[8]), .B(partialProduct_28[7]), .Cin(partialProduct_29[6]));
wire wire_592, wire_593;
bit_adder add277(.S(wire_592), .Cout(wire_593),  .A(partialProduct_27[9]), .B(partialProduct_28[8]), .Cin(partialProduct_29[7]));
wire wire_594, wire_595;
bit_adder add278(.S(wire_594), .Cout(wire_595),  .A(partialProduct_27[10]), .B(partialProduct_28[9]), .Cin(partialProduct_29[8]));
wire wire_596, wire_597;
bit_adder add279(.S(wire_596), .Cout(wire_597),  .A(partialProduct_27[11]), .B(partialProduct_28[10]), .Cin(partialProduct_29[9]));
wire wire_598, wire_599;
bit_adder add280(.S(wire_598), .Cout(wire_599),  .A(partialProduct_27[12]), .B(partialProduct_28[11]), .Cin(partialProduct_29[10]));
wire wire_600, wire_601;
bit_adder add281(.S(wire_600), .Cout(wire_601),  .A(partialProduct_27[13]), .B(partialProduct_28[12]), .Cin(partialProduct_29[11]));
wire wire_602, wire_603;
bit_adder add282(.S(wire_602), .Cout(wire_603),  .A(partialProduct_27[14]), .B(partialProduct_28[13]), .Cin(partialProduct_29[12]));
wire wire_604, wire_605;
bit_adder add283(.S(wire_604), .Cout(wire_605),  .A(partialProduct_27[15]), .B(partialProduct_28[14]), .Cin(partialProduct_29[13]));
wire wire_606, wire_607;
bit_adder add284(.S(wire_606), .Cout(wire_607),  .A(partialProduct_27[16]), .B(partialProduct_28[15]), .Cin(partialProduct_29[14]));
wire wire_608, wire_609;
bit_adder add285(.S(wire_608), .Cout(wire_609),  .A(partialProduct_27[17]), .B(partialProduct_28[16]), .Cin(partialProduct_29[15]));
wire wire_610, wire_611;
bit_adder add286(.S(wire_610), .Cout(wire_611),  .A(partialProduct_27[18]), .B(partialProduct_28[17]), .Cin(partialProduct_29[16]));
wire wire_612, wire_613;
bit_adder add287(.S(wire_612), .Cout(wire_613),  .A(partialProduct_27[19]), .B(partialProduct_28[18]), .Cin(partialProduct_29[17]));
wire wire_614, wire_615;
bit_adder add288(.S(wire_614), .Cout(wire_615),  .A(partialProduct_27[20]), .B(partialProduct_28[19]), .Cin(partialProduct_29[18]));
wire wire_616, wire_617;
bit_adder add289(.S(wire_616), .Cout(wire_617),  .A(partialProduct_27[21]), .B(partialProduct_28[20]), .Cin(partialProduct_29[19]));
wire wire_618, wire_619;
bit_adder add290(.S(wire_618), .Cout(wire_619),  .A(partialProduct_27[22]), .B(partialProduct_28[21]), .Cin(partialProduct_29[20]));
wire wire_620, wire_621;
bit_adder add291(.S(wire_620), .Cout(wire_621),  .A(partialProduct_27[23]), .B(partialProduct_28[22]), .Cin(partialProduct_29[21]));
wire wire_622, wire_623;
bit_adder add292(.S(wire_622), .Cout(wire_623),  .A(partialProduct_27[24]), .B(partialProduct_28[23]), .Cin(partialProduct_29[22]));
wire wire_624, wire_625;
bit_adder add293(.S(wire_624), .Cout(wire_625),  .A(partialProduct_27[25]), .B(partialProduct_28[24]), .Cin(partialProduct_29[23]));
wire wire_626, wire_627;
bit_adder add294(.S(wire_626), .Cout(wire_627),  .A(partialProduct_27[26]), .B(partialProduct_28[25]), .Cin(partialProduct_29[24]));
wire wire_628, wire_629;
bit_adder add295(.S(wire_628), .Cout(wire_629),  .A(partialProduct_27[27]), .B(partialProduct_28[26]), .Cin(partialProduct_29[25]));
wire wire_630, wire_631;
bit_adder add296(.S(wire_630), .Cout(wire_631),  .A(partialProduct_27[28]), .B(partialProduct_28[27]), .Cin(partialProduct_29[26]));
wire wire_632, wire_633;
bit_adder add297(.S(wire_632), .Cout(wire_633),  .A(partialProduct_27[29]), .B(partialProduct_28[28]), .Cin(partialProduct_29[27]));
wire wire_634, wire_635;
bit_adder add298(.S(wire_634), .Cout(wire_635),  .A(partialProduct_27[30]), .B(partialProduct_28[29]), .Cin(partialProduct_29[28]));
wire wire_636, wire_637;
bit_adder add299(.S(wire_636), .Cout(wire_637),  .A(partialProduct_27[31]), .B(partialProduct_28[30]), .Cin(partialProduct_29[29]));
wire wire_638, wire_639;
assign wire_638 = partialProduct_28[31] ^ partialProduct_29[30];
assign wire_639 = partialProduct_28[31] & partialProduct_29[30];
wire wire_640, wire_641;
assign wire_640 = wire_2 ^ wire_1;
assign wire_641 = wire_2 & wire_1;
wire wire_642, wire_643;
bit_adder add300(.S(wire_642), .Cout(wire_643),  .A(wire_4), .B(wire_3), .Cin(partialProduct_3[0]));
wire wire_644, wire_645;
bit_adder add301(.S(wire_644), .Cout(wire_645),  .A(wire_6), .B(wire_5), .Cin(wire_64));
wire wire_646, wire_647;
bit_adder add302(.S(wire_646), .Cout(wire_647),  .A(wire_8), .B(wire_7), .Cin(wire_66));
wire wire_648, wire_649;
bit_adder add303(.S(wire_648), .Cout(wire_649),  .A(wire_10), .B(wire_9), .Cin(wire_68));
wire wire_650, wire_651;
bit_adder add304(.S(wire_650), .Cout(wire_651),  .A(wire_12), .B(wire_11), .Cin(wire_70));
wire wire_652, wire_653;
bit_adder add305(.S(wire_652), .Cout(wire_653),  .A(wire_14), .B(wire_13), .Cin(wire_72));
wire wire_654, wire_655;
bit_adder add306(.S(wire_654), .Cout(wire_655),  .A(wire_16), .B(wire_15), .Cin(wire_74));
wire wire_656, wire_657;
bit_adder add307(.S(wire_656), .Cout(wire_657),  .A(wire_18), .B(wire_17), .Cin(wire_76));
wire wire_658, wire_659;
bit_adder add308(.S(wire_658), .Cout(wire_659),  .A(wire_20), .B(wire_19), .Cin(wire_78));
wire wire_660, wire_661;
bit_adder add309(.S(wire_660), .Cout(wire_661),  .A(wire_22), .B(wire_21), .Cin(wire_80));
wire wire_662, wire_663;
bit_adder add310(.S(wire_662), .Cout(wire_663),  .A(wire_24), .B(wire_23), .Cin(wire_82));
wire wire_664, wire_665;
bit_adder add311(.S(wire_664), .Cout(wire_665),  .A(wire_26), .B(wire_25), .Cin(wire_84));
wire wire_666, wire_667;
bit_adder add312(.S(wire_666), .Cout(wire_667),  .A(wire_28), .B(wire_27), .Cin(wire_86));
wire wire_668, wire_669;
bit_adder add313(.S(wire_668), .Cout(wire_669),  .A(wire_30), .B(wire_29), .Cin(wire_88));
wire wire_670, wire_671;
bit_adder add314(.S(wire_670), .Cout(wire_671),  .A(wire_32), .B(wire_31), .Cin(wire_90));
wire wire_672, wire_673;
bit_adder add315(.S(wire_672), .Cout(wire_673),  .A(wire_34), .B(wire_33), .Cin(wire_92));
wire wire_674, wire_675;
bit_adder add316(.S(wire_674), .Cout(wire_675),  .A(wire_36), .B(wire_35), .Cin(wire_94));
wire wire_676, wire_677;
bit_adder add317(.S(wire_676), .Cout(wire_677),  .A(wire_38), .B(wire_37), .Cin(wire_96));
wire wire_678, wire_679;
bit_adder add318(.S(wire_678), .Cout(wire_679),  .A(wire_40), .B(wire_39), .Cin(wire_98));
wire wire_680, wire_681;
bit_adder add319(.S(wire_680), .Cout(wire_681),  .A(wire_42), .B(wire_41), .Cin(wire_100));
wire wire_682, wire_683;
bit_adder add320(.S(wire_682), .Cout(wire_683),  .A(wire_44), .B(wire_43), .Cin(wire_102));
wire wire_684, wire_685;
bit_adder add321(.S(wire_684), .Cout(wire_685),  .A(wire_46), .B(wire_45), .Cin(wire_104));
wire wire_686, wire_687;
bit_adder add322(.S(wire_686), .Cout(wire_687),  .A(wire_48), .B(wire_47), .Cin(wire_106));
wire wire_688, wire_689;
bit_adder add323(.S(wire_688), .Cout(wire_689),  .A(wire_50), .B(wire_49), .Cin(wire_108));
wire wire_690, wire_691;
bit_adder add324(.S(wire_690), .Cout(wire_691),  .A(wire_52), .B(wire_51), .Cin(wire_110));
wire wire_692, wire_693;
bit_adder add325(.S(wire_692), .Cout(wire_693),  .A(wire_54), .B(wire_53), .Cin(wire_112));
wire wire_694, wire_695;
bit_adder add326(.S(wire_694), .Cout(wire_695),  .A(wire_56), .B(wire_55), .Cin(wire_114));
wire wire_696, wire_697;
bit_adder add327(.S(wire_696), .Cout(wire_697),  .A(wire_58), .B(wire_57), .Cin(wire_116));
wire wire_698, wire_699;
bit_adder add328(.S(wire_698), .Cout(wire_699),  .A(wire_60), .B(wire_59), .Cin(wire_118));
wire wire_700, wire_701;
bit_adder add329(.S(wire_700), .Cout(wire_701),  .A(wire_62), .B(wire_61), .Cin(wire_120));
wire wire_702, wire_703;
bit_adder add330(.S(wire_702), .Cout(wire_703),  .A(partialProduct_2[31]), .B(wire_63), .Cin(wire_122));
wire wire_704, wire_705;
assign wire_704 = wire_67 ^ partialProduct_6[0];
assign wire_705 = wire_67 & partialProduct_6[0];
wire wire_706, wire_707;
assign wire_706 = wire_69 ^ wire_128;
assign wire_707 = wire_69 & wire_128;
wire wire_708, wire_709;
bit_adder add331(.S(wire_708), .Cout(wire_709),  .A(wire_71), .B(wire_130), .Cin(wire_129));
wire wire_710, wire_711;
bit_adder add332(.S(wire_710), .Cout(wire_711),  .A(wire_73), .B(wire_132), .Cin(wire_131));
wire wire_712, wire_713;
bit_adder add333(.S(wire_712), .Cout(wire_713),  .A(wire_75), .B(wire_134), .Cin(wire_133));
wire wire_714, wire_715;
bit_adder add334(.S(wire_714), .Cout(wire_715),  .A(wire_77), .B(wire_136), .Cin(wire_135));
wire wire_716, wire_717;
bit_adder add335(.S(wire_716), .Cout(wire_717),  .A(wire_79), .B(wire_138), .Cin(wire_137));
wire wire_718, wire_719;
bit_adder add336(.S(wire_718), .Cout(wire_719),  .A(wire_81), .B(wire_140), .Cin(wire_139));
wire wire_720, wire_721;
bit_adder add337(.S(wire_720), .Cout(wire_721),  .A(wire_83), .B(wire_142), .Cin(wire_141));
wire wire_722, wire_723;
bit_adder add338(.S(wire_722), .Cout(wire_723),  .A(wire_85), .B(wire_144), .Cin(wire_143));
wire wire_724, wire_725;
bit_adder add339(.S(wire_724), .Cout(wire_725),  .A(wire_87), .B(wire_146), .Cin(wire_145));
wire wire_726, wire_727;
bit_adder add340(.S(wire_726), .Cout(wire_727),  .A(wire_89), .B(wire_148), .Cin(wire_147));
wire wire_728, wire_729;
bit_adder add341(.S(wire_728), .Cout(wire_729),  .A(wire_91), .B(wire_150), .Cin(wire_149));
wire wire_730, wire_731;
bit_adder add342(.S(wire_730), .Cout(wire_731),  .A(wire_93), .B(wire_152), .Cin(wire_151));
wire wire_732, wire_733;
bit_adder add343(.S(wire_732), .Cout(wire_733),  .A(wire_95), .B(wire_154), .Cin(wire_153));
wire wire_734, wire_735;
bit_adder add344(.S(wire_734), .Cout(wire_735),  .A(wire_97), .B(wire_156), .Cin(wire_155));
wire wire_736, wire_737;
bit_adder add345(.S(wire_736), .Cout(wire_737),  .A(wire_99), .B(wire_158), .Cin(wire_157));
wire wire_738, wire_739;
bit_adder add346(.S(wire_738), .Cout(wire_739),  .A(wire_101), .B(wire_160), .Cin(wire_159));
wire wire_740, wire_741;
bit_adder add347(.S(wire_740), .Cout(wire_741),  .A(wire_103), .B(wire_162), .Cin(wire_161));
wire wire_742, wire_743;
bit_adder add348(.S(wire_742), .Cout(wire_743),  .A(wire_105), .B(wire_164), .Cin(wire_163));
wire wire_744, wire_745;
bit_adder add349(.S(wire_744), .Cout(wire_745),  .A(wire_107), .B(wire_166), .Cin(wire_165));
wire wire_746, wire_747;
bit_adder add350(.S(wire_746), .Cout(wire_747),  .A(wire_109), .B(wire_168), .Cin(wire_167));
wire wire_748, wire_749;
bit_adder add351(.S(wire_748), .Cout(wire_749),  .A(wire_111), .B(wire_170), .Cin(wire_169));
wire wire_750, wire_751;
bit_adder add352(.S(wire_750), .Cout(wire_751),  .A(wire_113), .B(wire_172), .Cin(wire_171));
wire wire_752, wire_753;
bit_adder add353(.S(wire_752), .Cout(wire_753),  .A(wire_115), .B(wire_174), .Cin(wire_173));
wire wire_754, wire_755;
bit_adder add354(.S(wire_754), .Cout(wire_755),  .A(wire_117), .B(wire_176), .Cin(wire_175));
wire wire_756, wire_757;
bit_adder add355(.S(wire_756), .Cout(wire_757),  .A(wire_119), .B(wire_178), .Cin(wire_177));
wire wire_758, wire_759;
bit_adder add356(.S(wire_758), .Cout(wire_759),  .A(wire_121), .B(wire_180), .Cin(wire_179));
wire wire_760, wire_761;
bit_adder add357(.S(wire_760), .Cout(wire_761),  .A(wire_123), .B(wire_182), .Cin(wire_181));
wire wire_762, wire_763;
bit_adder add358(.S(wire_762), .Cout(wire_763),  .A(wire_125), .B(wire_184), .Cin(wire_183));
wire wire_764, wire_765;
bit_adder add359(.S(wire_764), .Cout(wire_765),  .A(wire_127), .B(wire_186), .Cin(wire_185));
wire wire_766, wire_767;
assign wire_766 = wire_188 ^ wire_187;
assign wire_767 = wire_188 & wire_187;
wire wire_768, wire_769;
assign wire_768 = wire_190 ^ wire_189;
assign wire_769 = wire_190 & wire_189;
wire wire_770, wire_771;
assign wire_770 = partialProduct_8[31] ^ wire_191;
assign wire_771 = partialProduct_8[31] & wire_191;
wire wire_772, wire_773;
assign wire_772 = wire_194 ^ wire_193;
assign wire_773 = wire_194 & wire_193;
wire wire_774, wire_775;
bit_adder add360(.S(wire_774), .Cout(wire_775),  .A(wire_196), .B(wire_195), .Cin(partialProduct_12[0]));
wire wire_776, wire_777;
bit_adder add361(.S(wire_776), .Cout(wire_777),  .A(wire_198), .B(wire_197), .Cin(wire_256));
wire wire_778, wire_779;
bit_adder add362(.S(wire_778), .Cout(wire_779),  .A(wire_200), .B(wire_199), .Cin(wire_258));
wire wire_780, wire_781;
bit_adder add363(.S(wire_780), .Cout(wire_781),  .A(wire_202), .B(wire_201), .Cin(wire_260));
wire wire_782, wire_783;
bit_adder add364(.S(wire_782), .Cout(wire_783),  .A(wire_204), .B(wire_203), .Cin(wire_262));
wire wire_784, wire_785;
bit_adder add365(.S(wire_784), .Cout(wire_785),  .A(wire_206), .B(wire_205), .Cin(wire_264));
wire wire_786, wire_787;
bit_adder add366(.S(wire_786), .Cout(wire_787),  .A(wire_208), .B(wire_207), .Cin(wire_266));
wire wire_788, wire_789;
bit_adder add367(.S(wire_788), .Cout(wire_789),  .A(wire_210), .B(wire_209), .Cin(wire_268));
wire wire_790, wire_791;
bit_adder add368(.S(wire_790), .Cout(wire_791),  .A(wire_212), .B(wire_211), .Cin(wire_270));
wire wire_792, wire_793;
bit_adder add369(.S(wire_792), .Cout(wire_793),  .A(wire_214), .B(wire_213), .Cin(wire_272));
wire wire_794, wire_795;
bit_adder add370(.S(wire_794), .Cout(wire_795),  .A(wire_216), .B(wire_215), .Cin(wire_274));
wire wire_796, wire_797;
bit_adder add371(.S(wire_796), .Cout(wire_797),  .A(wire_218), .B(wire_217), .Cin(wire_276));
wire wire_798, wire_799;
bit_adder add372(.S(wire_798), .Cout(wire_799),  .A(wire_220), .B(wire_219), .Cin(wire_278));
wire wire_800, wire_801;
bit_adder add373(.S(wire_800), .Cout(wire_801),  .A(wire_222), .B(wire_221), .Cin(wire_280));
wire wire_802, wire_803;
bit_adder add374(.S(wire_802), .Cout(wire_803),  .A(wire_224), .B(wire_223), .Cin(wire_282));
wire wire_804, wire_805;
bit_adder add375(.S(wire_804), .Cout(wire_805),  .A(wire_226), .B(wire_225), .Cin(wire_284));
wire wire_806, wire_807;
bit_adder add376(.S(wire_806), .Cout(wire_807),  .A(wire_228), .B(wire_227), .Cin(wire_286));
wire wire_808, wire_809;
bit_adder add377(.S(wire_808), .Cout(wire_809),  .A(wire_230), .B(wire_229), .Cin(wire_288));
wire wire_810, wire_811;
bit_adder add378(.S(wire_810), .Cout(wire_811),  .A(wire_232), .B(wire_231), .Cin(wire_290));
wire wire_812, wire_813;
bit_adder add379(.S(wire_812), .Cout(wire_813),  .A(wire_234), .B(wire_233), .Cin(wire_292));
wire wire_814, wire_815;
bit_adder add380(.S(wire_814), .Cout(wire_815),  .A(wire_236), .B(wire_235), .Cin(wire_294));
wire wire_816, wire_817;
bit_adder add381(.S(wire_816), .Cout(wire_817),  .A(wire_238), .B(wire_237), .Cin(wire_296));
wire wire_818, wire_819;
bit_adder add382(.S(wire_818), .Cout(wire_819),  .A(wire_240), .B(wire_239), .Cin(wire_298));
wire wire_820, wire_821;
bit_adder add383(.S(wire_820), .Cout(wire_821),  .A(wire_242), .B(wire_241), .Cin(wire_300));
wire wire_822, wire_823;
bit_adder add384(.S(wire_822), .Cout(wire_823),  .A(wire_244), .B(wire_243), .Cin(wire_302));
wire wire_824, wire_825;
bit_adder add385(.S(wire_824), .Cout(wire_825),  .A(wire_246), .B(wire_245), .Cin(wire_304));
wire wire_826, wire_827;
bit_adder add386(.S(wire_826), .Cout(wire_827),  .A(wire_248), .B(wire_247), .Cin(wire_306));
wire wire_828, wire_829;
bit_adder add387(.S(wire_828), .Cout(wire_829),  .A(wire_250), .B(wire_249), .Cin(wire_308));
wire wire_830, wire_831;
bit_adder add388(.S(wire_830), .Cout(wire_831),  .A(wire_252), .B(wire_251), .Cin(wire_310));
wire wire_832, wire_833;
bit_adder add389(.S(wire_832), .Cout(wire_833),  .A(wire_254), .B(wire_253), .Cin(wire_312));
wire wire_834, wire_835;
bit_adder add390(.S(wire_834), .Cout(wire_835),  .A(partialProduct_11[31]), .B(wire_255), .Cin(wire_314));
wire wire_836, wire_837;
assign wire_836 = wire_259 ^ partialProduct_15[0];
assign wire_837 = wire_259 & partialProduct_15[0];
wire wire_838, wire_839;
assign wire_838 = wire_261 ^ wire_320;
assign wire_839 = wire_261 & wire_320;
wire wire_840, wire_841;
bit_adder add391(.S(wire_840), .Cout(wire_841),  .A(wire_263), .B(wire_322), .Cin(wire_321));
wire wire_842, wire_843;
bit_adder add392(.S(wire_842), .Cout(wire_843),  .A(wire_265), .B(wire_324), .Cin(wire_323));
wire wire_844, wire_845;
bit_adder add393(.S(wire_844), .Cout(wire_845),  .A(wire_267), .B(wire_326), .Cin(wire_325));
wire wire_846, wire_847;
bit_adder add394(.S(wire_846), .Cout(wire_847),  .A(wire_269), .B(wire_328), .Cin(wire_327));
wire wire_848, wire_849;
bit_adder add395(.S(wire_848), .Cout(wire_849),  .A(wire_271), .B(wire_330), .Cin(wire_329));
wire wire_850, wire_851;
bit_adder add396(.S(wire_850), .Cout(wire_851),  .A(wire_273), .B(wire_332), .Cin(wire_331));
wire wire_852, wire_853;
bit_adder add397(.S(wire_852), .Cout(wire_853),  .A(wire_275), .B(wire_334), .Cin(wire_333));
wire wire_854, wire_855;
bit_adder add398(.S(wire_854), .Cout(wire_855),  .A(wire_277), .B(wire_336), .Cin(wire_335));
wire wire_856, wire_857;
bit_adder add399(.S(wire_856), .Cout(wire_857),  .A(wire_279), .B(wire_338), .Cin(wire_337));
wire wire_858, wire_859;
bit_adder add400(.S(wire_858), .Cout(wire_859),  .A(wire_281), .B(wire_340), .Cin(wire_339));
wire wire_860, wire_861;
bit_adder add401(.S(wire_860), .Cout(wire_861),  .A(wire_283), .B(wire_342), .Cin(wire_341));
wire wire_862, wire_863;
bit_adder add402(.S(wire_862), .Cout(wire_863),  .A(wire_285), .B(wire_344), .Cin(wire_343));
wire wire_864, wire_865;
bit_adder add403(.S(wire_864), .Cout(wire_865),  .A(wire_287), .B(wire_346), .Cin(wire_345));
wire wire_866, wire_867;
bit_adder add404(.S(wire_866), .Cout(wire_867),  .A(wire_289), .B(wire_348), .Cin(wire_347));
wire wire_868, wire_869;
bit_adder add405(.S(wire_868), .Cout(wire_869),  .A(wire_291), .B(wire_350), .Cin(wire_349));
wire wire_870, wire_871;
bit_adder add406(.S(wire_870), .Cout(wire_871),  .A(wire_293), .B(wire_352), .Cin(wire_351));
wire wire_872, wire_873;
bit_adder add407(.S(wire_872), .Cout(wire_873),  .A(wire_295), .B(wire_354), .Cin(wire_353));
wire wire_874, wire_875;
bit_adder add408(.S(wire_874), .Cout(wire_875),  .A(wire_297), .B(wire_356), .Cin(wire_355));
wire wire_876, wire_877;
bit_adder add409(.S(wire_876), .Cout(wire_877),  .A(wire_299), .B(wire_358), .Cin(wire_357));
wire wire_878, wire_879;
bit_adder add410(.S(wire_878), .Cout(wire_879),  .A(wire_301), .B(wire_360), .Cin(wire_359));
wire wire_880, wire_881;
bit_adder add411(.S(wire_880), .Cout(wire_881),  .A(wire_303), .B(wire_362), .Cin(wire_361));
wire wire_882, wire_883;
bit_adder add412(.S(wire_882), .Cout(wire_883),  .A(wire_305), .B(wire_364), .Cin(wire_363));
wire wire_884, wire_885;
bit_adder add413(.S(wire_884), .Cout(wire_885),  .A(wire_307), .B(wire_366), .Cin(wire_365));
wire wire_886, wire_887;
bit_adder add414(.S(wire_886), .Cout(wire_887),  .A(wire_309), .B(wire_368), .Cin(wire_367));
wire wire_888, wire_889;
bit_adder add415(.S(wire_888), .Cout(wire_889),  .A(wire_311), .B(wire_370), .Cin(wire_369));
wire wire_890, wire_891;
bit_adder add416(.S(wire_890), .Cout(wire_891),  .A(wire_313), .B(wire_372), .Cin(wire_371));
wire wire_892, wire_893;
bit_adder add417(.S(wire_892), .Cout(wire_893),  .A(wire_315), .B(wire_374), .Cin(wire_373));
wire wire_894, wire_895;
bit_adder add418(.S(wire_894), .Cout(wire_895),  .A(wire_317), .B(wire_376), .Cin(wire_375));
wire wire_896, wire_897;
bit_adder add419(.S(wire_896), .Cout(wire_897),  .A(wire_319), .B(wire_378), .Cin(wire_377));
wire wire_898, wire_899;
assign wire_898 = wire_380 ^ wire_379;
assign wire_899 = wire_380 & wire_379;
wire wire_900, wire_901;
assign wire_900 = wire_382 ^ wire_381;
assign wire_901 = wire_382 & wire_381;
wire wire_902, wire_903;
assign wire_902 = partialProduct_17[31] ^ wire_383;
assign wire_903 = partialProduct_17[31] & wire_383;
wire wire_904, wire_905;
assign wire_904 = wire_386 ^ wire_385;
assign wire_905 = wire_386 & wire_385;
wire wire_906, wire_907;
bit_adder add420(.S(wire_906), .Cout(wire_907),  .A(wire_388), .B(wire_387), .Cin(partialProduct_21[0]));
wire wire_908, wire_909;
bit_adder add421(.S(wire_908), .Cout(wire_909),  .A(wire_390), .B(wire_389), .Cin(wire_448));
wire wire_910, wire_911;
bit_adder add422(.S(wire_910), .Cout(wire_911),  .A(wire_392), .B(wire_391), .Cin(wire_450));
wire wire_912, wire_913;
bit_adder add423(.S(wire_912), .Cout(wire_913),  .A(wire_394), .B(wire_393), .Cin(wire_452));
wire wire_914, wire_915;
bit_adder add424(.S(wire_914), .Cout(wire_915),  .A(wire_396), .B(wire_395), .Cin(wire_454));
wire wire_916, wire_917;
bit_adder add425(.S(wire_916), .Cout(wire_917),  .A(wire_398), .B(wire_397), .Cin(wire_456));
wire wire_918, wire_919;
bit_adder add426(.S(wire_918), .Cout(wire_919),  .A(wire_400), .B(wire_399), .Cin(wire_458));
wire wire_920, wire_921;
bit_adder add427(.S(wire_920), .Cout(wire_921),  .A(wire_402), .B(wire_401), .Cin(wire_460));
wire wire_922, wire_923;
bit_adder add428(.S(wire_922), .Cout(wire_923),  .A(wire_404), .B(wire_403), .Cin(wire_462));
wire wire_924, wire_925;
bit_adder add429(.S(wire_924), .Cout(wire_925),  .A(wire_406), .B(wire_405), .Cin(wire_464));
wire wire_926, wire_927;
bit_adder add430(.S(wire_926), .Cout(wire_927),  .A(wire_408), .B(wire_407), .Cin(wire_466));
wire wire_928, wire_929;
bit_adder add431(.S(wire_928), .Cout(wire_929),  .A(wire_410), .B(wire_409), .Cin(wire_468));
wire wire_930, wire_931;
bit_adder add432(.S(wire_930), .Cout(wire_931),  .A(wire_412), .B(wire_411), .Cin(wire_470));
wire wire_932, wire_933;
bit_adder add433(.S(wire_932), .Cout(wire_933),  .A(wire_414), .B(wire_413), .Cin(wire_472));
wire wire_934, wire_935;
bit_adder add434(.S(wire_934), .Cout(wire_935),  .A(wire_416), .B(wire_415), .Cin(wire_474));
wire wire_936, wire_937;
bit_adder add435(.S(wire_936), .Cout(wire_937),  .A(wire_418), .B(wire_417), .Cin(wire_476));
wire wire_938, wire_939;
bit_adder add436(.S(wire_938), .Cout(wire_939),  .A(wire_420), .B(wire_419), .Cin(wire_478));
wire wire_940, wire_941;
bit_adder add437(.S(wire_940), .Cout(wire_941),  .A(wire_422), .B(wire_421), .Cin(wire_480));
wire wire_942, wire_943;
bit_adder add438(.S(wire_942), .Cout(wire_943),  .A(wire_424), .B(wire_423), .Cin(wire_482));
wire wire_944, wire_945;
bit_adder add439(.S(wire_944), .Cout(wire_945),  .A(wire_426), .B(wire_425), .Cin(wire_484));
wire wire_946, wire_947;
bit_adder add440(.S(wire_946), .Cout(wire_947),  .A(wire_428), .B(wire_427), .Cin(wire_486));
wire wire_948, wire_949;
bit_adder add441(.S(wire_948), .Cout(wire_949),  .A(wire_430), .B(wire_429), .Cin(wire_488));
wire wire_950, wire_951;
bit_adder add442(.S(wire_950), .Cout(wire_951),  .A(wire_432), .B(wire_431), .Cin(wire_490));
wire wire_952, wire_953;
bit_adder add443(.S(wire_952), .Cout(wire_953),  .A(wire_434), .B(wire_433), .Cin(wire_492));
wire wire_954, wire_955;
bit_adder add444(.S(wire_954), .Cout(wire_955),  .A(wire_436), .B(wire_435), .Cin(wire_494));
wire wire_956, wire_957;
bit_adder add445(.S(wire_956), .Cout(wire_957),  .A(wire_438), .B(wire_437), .Cin(wire_496));
wire wire_958, wire_959;
bit_adder add446(.S(wire_958), .Cout(wire_959),  .A(wire_440), .B(wire_439), .Cin(wire_498));
wire wire_960, wire_961;
bit_adder add447(.S(wire_960), .Cout(wire_961),  .A(wire_442), .B(wire_441), .Cin(wire_500));
wire wire_962, wire_963;
bit_adder add448(.S(wire_962), .Cout(wire_963),  .A(wire_444), .B(wire_443), .Cin(wire_502));
wire wire_964, wire_965;
bit_adder add449(.S(wire_964), .Cout(wire_965),  .A(wire_446), .B(wire_445), .Cin(wire_504));
wire wire_966, wire_967;
bit_adder add450(.S(wire_966), .Cout(wire_967),  .A(partialProduct_20[31]), .B(wire_447), .Cin(wire_506));
wire wire_968, wire_969;
assign wire_968 = wire_451 ^ partialProduct_24[0];
assign wire_969 = wire_451 & partialProduct_24[0];
wire wire_970, wire_971;
assign wire_970 = wire_453 ^ wire_512;
assign wire_971 = wire_453 & wire_512;
wire wire_972, wire_973;
bit_adder add451(.S(wire_972), .Cout(wire_973),  .A(wire_455), .B(wire_514), .Cin(wire_513));
wire wire_974, wire_975;
bit_adder add452(.S(wire_974), .Cout(wire_975),  .A(wire_457), .B(wire_516), .Cin(wire_515));
wire wire_976, wire_977;
bit_adder add453(.S(wire_976), .Cout(wire_977),  .A(wire_459), .B(wire_518), .Cin(wire_517));
wire wire_978, wire_979;
bit_adder add454(.S(wire_978), .Cout(wire_979),  .A(wire_461), .B(wire_520), .Cin(wire_519));
wire wire_980, wire_981;
bit_adder add455(.S(wire_980), .Cout(wire_981),  .A(wire_463), .B(wire_522), .Cin(wire_521));
wire wire_982, wire_983;
bit_adder add456(.S(wire_982), .Cout(wire_983),  .A(wire_465), .B(wire_524), .Cin(wire_523));
wire wire_984, wire_985;
bit_adder add457(.S(wire_984), .Cout(wire_985),  .A(wire_467), .B(wire_526), .Cin(wire_525));
wire wire_986, wire_987;
bit_adder add458(.S(wire_986), .Cout(wire_987),  .A(wire_469), .B(wire_528), .Cin(wire_527));
wire wire_988, wire_989;
bit_adder add459(.S(wire_988), .Cout(wire_989),  .A(wire_471), .B(wire_530), .Cin(wire_529));
wire wire_990, wire_991;
bit_adder add460(.S(wire_990), .Cout(wire_991),  .A(wire_473), .B(wire_532), .Cin(wire_531));
wire wire_992, wire_993;
bit_adder add461(.S(wire_992), .Cout(wire_993),  .A(wire_475), .B(wire_534), .Cin(wire_533));
wire wire_994, wire_995;
bit_adder add462(.S(wire_994), .Cout(wire_995),  .A(wire_477), .B(wire_536), .Cin(wire_535));
wire wire_996, wire_997;
bit_adder add463(.S(wire_996), .Cout(wire_997),  .A(wire_479), .B(wire_538), .Cin(wire_537));
wire wire_998, wire_999;
bit_adder add464(.S(wire_998), .Cout(wire_999),  .A(wire_481), .B(wire_540), .Cin(wire_539));
wire wire_1000, wire_1001;
bit_adder add465(.S(wire_1000), .Cout(wire_1001),  .A(wire_483), .B(wire_542), .Cin(wire_541));
wire wire_1002, wire_1003;
bit_adder add466(.S(wire_1002), .Cout(wire_1003),  .A(wire_485), .B(wire_544), .Cin(wire_543));
wire wire_1004, wire_1005;
bit_adder add467(.S(wire_1004), .Cout(wire_1005),  .A(wire_487), .B(wire_546), .Cin(wire_545));
wire wire_1006, wire_1007;
bit_adder add468(.S(wire_1006), .Cout(wire_1007),  .A(wire_489), .B(wire_548), .Cin(wire_547));
wire wire_1008, wire_1009;
bit_adder add469(.S(wire_1008), .Cout(wire_1009),  .A(wire_491), .B(wire_550), .Cin(wire_549));
wire wire_1010, wire_1011;
bit_adder add470(.S(wire_1010), .Cout(wire_1011),  .A(wire_493), .B(wire_552), .Cin(wire_551));
wire wire_1012, wire_1013;
bit_adder add471(.S(wire_1012), .Cout(wire_1013),  .A(wire_495), .B(wire_554), .Cin(wire_553));
wire wire_1014, wire_1015;
bit_adder add472(.S(wire_1014), .Cout(wire_1015),  .A(wire_497), .B(wire_556), .Cin(wire_555));
wire wire_1016, wire_1017;
bit_adder add473(.S(wire_1016), .Cout(wire_1017),  .A(wire_499), .B(wire_558), .Cin(wire_557));
wire wire_1018, wire_1019;
bit_adder add474(.S(wire_1018), .Cout(wire_1019),  .A(wire_501), .B(wire_560), .Cin(wire_559));
wire wire_1020, wire_1021;
bit_adder add475(.S(wire_1020), .Cout(wire_1021),  .A(wire_503), .B(wire_562), .Cin(wire_561));
wire wire_1022, wire_1023;
bit_adder add476(.S(wire_1022), .Cout(wire_1023),  .A(wire_505), .B(wire_564), .Cin(wire_563));
wire wire_1024, wire_1025;
bit_adder add477(.S(wire_1024), .Cout(wire_1025),  .A(wire_507), .B(wire_566), .Cin(wire_565));
wire wire_1026, wire_1027;
bit_adder add478(.S(wire_1026), .Cout(wire_1027),  .A(wire_509), .B(wire_568), .Cin(wire_567));
wire wire_1028, wire_1029;
bit_adder add479(.S(wire_1028), .Cout(wire_1029),  .A(wire_511), .B(wire_570), .Cin(wire_569));
wire wire_1030, wire_1031;
assign wire_1030 = wire_572 ^ wire_571;
assign wire_1031 = wire_572 & wire_571;
wire wire_1032, wire_1033;
assign wire_1032 = wire_574 ^ wire_573;
assign wire_1033 = wire_574 & wire_573;
wire wire_1034, wire_1035;
assign wire_1034 = partialProduct_26[31] ^ wire_575;
assign wire_1035 = partialProduct_26[31] & wire_575;
wire wire_1036, wire_1037;
assign wire_1036 = wire_578 ^ wire_577;
assign wire_1037 = wire_578 & wire_577;
wire wire_1038, wire_1039;
bit_adder add480(.S(wire_1038), .Cout(wire_1039),  .A(wire_580), .B(wire_579), .Cin(partialProduct_30[0]));
wire wire_1040, wire_1041;
bit_adder add481(.S(wire_1040), .Cout(wire_1041),  .A(wire_582), .B(wire_581), .Cin(partialProduct_30[1]));
wire wire_1042, wire_1043;
bit_adder add482(.S(wire_1042), .Cout(wire_1043),  .A(wire_584), .B(wire_583), .Cin(partialProduct_30[2]));
wire wire_1044, wire_1045;
bit_adder add483(.S(wire_1044), .Cout(wire_1045),  .A(wire_586), .B(wire_585), .Cin(partialProduct_30[3]));
wire wire_1046, wire_1047;
bit_adder add484(.S(wire_1046), .Cout(wire_1047),  .A(wire_588), .B(wire_587), .Cin(partialProduct_30[4]));
wire wire_1048, wire_1049;
bit_adder add485(.S(wire_1048), .Cout(wire_1049),  .A(wire_590), .B(wire_589), .Cin(partialProduct_30[5]));
wire wire_1050, wire_1051;
bit_adder add486(.S(wire_1050), .Cout(wire_1051),  .A(wire_592), .B(wire_591), .Cin(partialProduct_30[6]));
wire wire_1052, wire_1053;
bit_adder add487(.S(wire_1052), .Cout(wire_1053),  .A(wire_594), .B(wire_593), .Cin(partialProduct_30[7]));
wire wire_1054, wire_1055;
bit_adder add488(.S(wire_1054), .Cout(wire_1055),  .A(wire_596), .B(wire_595), .Cin(partialProduct_30[8]));
wire wire_1056, wire_1057;
bit_adder add489(.S(wire_1056), .Cout(wire_1057),  .A(wire_598), .B(wire_597), .Cin(partialProduct_30[9]));
wire wire_1058, wire_1059;
bit_adder add490(.S(wire_1058), .Cout(wire_1059),  .A(wire_600), .B(wire_599), .Cin(partialProduct_30[10]));
wire wire_1060, wire_1061;
bit_adder add491(.S(wire_1060), .Cout(wire_1061),  .A(wire_602), .B(wire_601), .Cin(partialProduct_30[11]));
wire wire_1062, wire_1063;
bit_adder add492(.S(wire_1062), .Cout(wire_1063),  .A(wire_604), .B(wire_603), .Cin(partialProduct_30[12]));
wire wire_1064, wire_1065;
bit_adder add493(.S(wire_1064), .Cout(wire_1065),  .A(wire_606), .B(wire_605), .Cin(partialProduct_30[13]));
wire wire_1066, wire_1067;
bit_adder add494(.S(wire_1066), .Cout(wire_1067),  .A(wire_608), .B(wire_607), .Cin(partialProduct_30[14]));
wire wire_1068, wire_1069;
bit_adder add495(.S(wire_1068), .Cout(wire_1069),  .A(wire_610), .B(wire_609), .Cin(partialProduct_30[15]));
wire wire_1070, wire_1071;
bit_adder add496(.S(wire_1070), .Cout(wire_1071),  .A(wire_612), .B(wire_611), .Cin(partialProduct_30[16]));
wire wire_1072, wire_1073;
bit_adder add497(.S(wire_1072), .Cout(wire_1073),  .A(wire_614), .B(wire_613), .Cin(partialProduct_30[17]));
wire wire_1074, wire_1075;
bit_adder add498(.S(wire_1074), .Cout(wire_1075),  .A(wire_616), .B(wire_615), .Cin(partialProduct_30[18]));
wire wire_1076, wire_1077;
bit_adder add499(.S(wire_1076), .Cout(wire_1077),  .A(wire_618), .B(wire_617), .Cin(partialProduct_30[19]));
wire wire_1078, wire_1079;
bit_adder add500(.S(wire_1078), .Cout(wire_1079),  .A(wire_620), .B(wire_619), .Cin(partialProduct_30[20]));
wire wire_1080, wire_1081;
bit_adder add501(.S(wire_1080), .Cout(wire_1081),  .A(wire_622), .B(wire_621), .Cin(partialProduct_30[21]));
wire wire_1082, wire_1083;
bit_adder add502(.S(wire_1082), .Cout(wire_1083),  .A(wire_624), .B(wire_623), .Cin(partialProduct_30[22]));
wire wire_1084, wire_1085;
bit_adder add503(.S(wire_1084), .Cout(wire_1085),  .A(wire_626), .B(wire_625), .Cin(partialProduct_30[23]));
wire wire_1086, wire_1087;
bit_adder add504(.S(wire_1086), .Cout(wire_1087),  .A(wire_628), .B(wire_627), .Cin(partialProduct_30[24]));
wire wire_1088, wire_1089;
bit_adder add505(.S(wire_1088), .Cout(wire_1089),  .A(wire_630), .B(wire_629), .Cin(partialProduct_30[25]));
wire wire_1090, wire_1091;
bit_adder add506(.S(wire_1090), .Cout(wire_1091),  .A(wire_632), .B(wire_631), .Cin(partialProduct_30[26]));
wire wire_1092, wire_1093;
bit_adder add507(.S(wire_1092), .Cout(wire_1093),  .A(wire_634), .B(wire_633), .Cin(partialProduct_30[27]));
wire wire_1094, wire_1095;
bit_adder add508(.S(wire_1094), .Cout(wire_1095),  .A(wire_636), .B(wire_635), .Cin(partialProduct_30[28]));
wire wire_1096, wire_1097;
bit_adder add509(.S(wire_1096), .Cout(wire_1097),  .A(wire_638), .B(wire_637), .Cin(partialProduct_30[29]));
wire wire_1098, wire_1099;
bit_adder add510(.S(wire_1098), .Cout(wire_1099),  .A(partialProduct_29[31]), .B(wire_639), .Cin(partialProduct_30[30]));
wire wire_1100, wire_1101;
assign wire_1100 = wire_642 ^ wire_641;
assign wire_1101 = wire_642 & wire_641;
wire wire_1102, wire_1103;
assign wire_1102 = wire_644 ^ wire_643;
assign wire_1103 = wire_644 & wire_643;
wire wire_1104, wire_1105;
bit_adder add511(.S(wire_1104), .Cout(wire_1105),  .A(wire_646), .B(wire_645), .Cin(wire_65));
wire wire_1106, wire_1107;
bit_adder add512(.S(wire_1106), .Cout(wire_1107),  .A(wire_648), .B(wire_647), .Cin(wire_704));
wire wire_1108, wire_1109;
bit_adder add513(.S(wire_1108), .Cout(wire_1109),  .A(wire_650), .B(wire_649), .Cin(wire_706));
wire wire_1110, wire_1111;
bit_adder add514(.S(wire_1110), .Cout(wire_1111),  .A(wire_652), .B(wire_651), .Cin(wire_708));
wire wire_1112, wire_1113;
bit_adder add515(.S(wire_1112), .Cout(wire_1113),  .A(wire_654), .B(wire_653), .Cin(wire_710));
wire wire_1114, wire_1115;
bit_adder add516(.S(wire_1114), .Cout(wire_1115),  .A(wire_656), .B(wire_655), .Cin(wire_712));
wire wire_1116, wire_1117;
bit_adder add517(.S(wire_1116), .Cout(wire_1117),  .A(wire_658), .B(wire_657), .Cin(wire_714));
wire wire_1118, wire_1119;
bit_adder add518(.S(wire_1118), .Cout(wire_1119),  .A(wire_660), .B(wire_659), .Cin(wire_716));
wire wire_1120, wire_1121;
bit_adder add519(.S(wire_1120), .Cout(wire_1121),  .A(wire_662), .B(wire_661), .Cin(wire_718));
wire wire_1122, wire_1123;
bit_adder add520(.S(wire_1122), .Cout(wire_1123),  .A(wire_664), .B(wire_663), .Cin(wire_720));
wire wire_1124, wire_1125;
bit_adder add521(.S(wire_1124), .Cout(wire_1125),  .A(wire_666), .B(wire_665), .Cin(wire_722));
wire wire_1126, wire_1127;
bit_adder add522(.S(wire_1126), .Cout(wire_1127),  .A(wire_668), .B(wire_667), .Cin(wire_724));
wire wire_1128, wire_1129;
bit_adder add523(.S(wire_1128), .Cout(wire_1129),  .A(wire_670), .B(wire_669), .Cin(wire_726));
wire wire_1130, wire_1131;
bit_adder add524(.S(wire_1130), .Cout(wire_1131),  .A(wire_672), .B(wire_671), .Cin(wire_728));
wire wire_1132, wire_1133;
bit_adder add525(.S(wire_1132), .Cout(wire_1133),  .A(wire_674), .B(wire_673), .Cin(wire_730));
wire wire_1134, wire_1135;
bit_adder add526(.S(wire_1134), .Cout(wire_1135),  .A(wire_676), .B(wire_675), .Cin(wire_732));
wire wire_1136, wire_1137;
bit_adder add527(.S(wire_1136), .Cout(wire_1137),  .A(wire_678), .B(wire_677), .Cin(wire_734));
wire wire_1138, wire_1139;
bit_adder add528(.S(wire_1138), .Cout(wire_1139),  .A(wire_680), .B(wire_679), .Cin(wire_736));
wire wire_1140, wire_1141;
bit_adder add529(.S(wire_1140), .Cout(wire_1141),  .A(wire_682), .B(wire_681), .Cin(wire_738));
wire wire_1142, wire_1143;
bit_adder add530(.S(wire_1142), .Cout(wire_1143),  .A(wire_684), .B(wire_683), .Cin(wire_740));
wire wire_1144, wire_1145;
bit_adder add531(.S(wire_1144), .Cout(wire_1145),  .A(wire_686), .B(wire_685), .Cin(wire_742));
wire wire_1146, wire_1147;
bit_adder add532(.S(wire_1146), .Cout(wire_1147),  .A(wire_688), .B(wire_687), .Cin(wire_744));
wire wire_1148, wire_1149;
bit_adder add533(.S(wire_1148), .Cout(wire_1149),  .A(wire_690), .B(wire_689), .Cin(wire_746));
wire wire_1150, wire_1151;
bit_adder add534(.S(wire_1150), .Cout(wire_1151),  .A(wire_692), .B(wire_691), .Cin(wire_748));
wire wire_1152, wire_1153;
bit_adder add535(.S(wire_1152), .Cout(wire_1153),  .A(wire_694), .B(wire_693), .Cin(wire_750));
wire wire_1154, wire_1155;
bit_adder add536(.S(wire_1154), .Cout(wire_1155),  .A(wire_696), .B(wire_695), .Cin(wire_752));
wire wire_1156, wire_1157;
bit_adder add537(.S(wire_1156), .Cout(wire_1157),  .A(wire_698), .B(wire_697), .Cin(wire_754));
wire wire_1158, wire_1159;
bit_adder add538(.S(wire_1158), .Cout(wire_1159),  .A(wire_700), .B(wire_699), .Cin(wire_756));
wire wire_1160, wire_1161;
bit_adder add539(.S(wire_1160), .Cout(wire_1161),  .A(wire_702), .B(wire_701), .Cin(wire_758));
wire wire_1162, wire_1163;
bit_adder add540(.S(wire_1162), .Cout(wire_1163),  .A(wire_124), .B(wire_703), .Cin(wire_760));
wire wire_1164, wire_1165;
assign wire_1164 = wire_126 ^ wire_762;
assign wire_1165 = wire_126 & wire_762;
wire wire_1166, wire_1167;
assign wire_1166 = partialProduct_5[31] ^ wire_764;
assign wire_1167 = partialProduct_5[31] & wire_764;
wire wire_1168, wire_1169;
assign wire_1168 = wire_709 ^ partialProduct_9[0];
assign wire_1169 = wire_709 & partialProduct_9[0];
wire wire_1170, wire_1171;
assign wire_1170 = wire_711 ^ wire_192;
assign wire_1171 = wire_711 & wire_192;
wire wire_1172, wire_1173;
assign wire_1172 = wire_713 ^ wire_772;
assign wire_1173 = wire_713 & wire_772;
wire wire_1174, wire_1175;
bit_adder add541(.S(wire_1174), .Cout(wire_1175),  .A(wire_715), .B(wire_774), .Cin(wire_773));
wire wire_1176, wire_1177;
bit_adder add542(.S(wire_1176), .Cout(wire_1177),  .A(wire_717), .B(wire_776), .Cin(wire_775));
wire wire_1178, wire_1179;
bit_adder add543(.S(wire_1178), .Cout(wire_1179),  .A(wire_719), .B(wire_778), .Cin(wire_777));
wire wire_1180, wire_1181;
bit_adder add544(.S(wire_1180), .Cout(wire_1181),  .A(wire_721), .B(wire_780), .Cin(wire_779));
wire wire_1182, wire_1183;
bit_adder add545(.S(wire_1182), .Cout(wire_1183),  .A(wire_723), .B(wire_782), .Cin(wire_781));
wire wire_1184, wire_1185;
bit_adder add546(.S(wire_1184), .Cout(wire_1185),  .A(wire_725), .B(wire_784), .Cin(wire_783));
wire wire_1186, wire_1187;
bit_adder add547(.S(wire_1186), .Cout(wire_1187),  .A(wire_727), .B(wire_786), .Cin(wire_785));
wire wire_1188, wire_1189;
bit_adder add548(.S(wire_1188), .Cout(wire_1189),  .A(wire_729), .B(wire_788), .Cin(wire_787));
wire wire_1190, wire_1191;
bit_adder add549(.S(wire_1190), .Cout(wire_1191),  .A(wire_731), .B(wire_790), .Cin(wire_789));
wire wire_1192, wire_1193;
bit_adder add550(.S(wire_1192), .Cout(wire_1193),  .A(wire_733), .B(wire_792), .Cin(wire_791));
wire wire_1194, wire_1195;
bit_adder add551(.S(wire_1194), .Cout(wire_1195),  .A(wire_735), .B(wire_794), .Cin(wire_793));
wire wire_1196, wire_1197;
bit_adder add552(.S(wire_1196), .Cout(wire_1197),  .A(wire_737), .B(wire_796), .Cin(wire_795));
wire wire_1198, wire_1199;
bit_adder add553(.S(wire_1198), .Cout(wire_1199),  .A(wire_739), .B(wire_798), .Cin(wire_797));
wire wire_1200, wire_1201;
bit_adder add554(.S(wire_1200), .Cout(wire_1201),  .A(wire_741), .B(wire_800), .Cin(wire_799));
wire wire_1202, wire_1203;
bit_adder add555(.S(wire_1202), .Cout(wire_1203),  .A(wire_743), .B(wire_802), .Cin(wire_801));
wire wire_1204, wire_1205;
bit_adder add556(.S(wire_1204), .Cout(wire_1205),  .A(wire_745), .B(wire_804), .Cin(wire_803));
wire wire_1206, wire_1207;
bit_adder add557(.S(wire_1206), .Cout(wire_1207),  .A(wire_747), .B(wire_806), .Cin(wire_805));
wire wire_1208, wire_1209;
bit_adder add558(.S(wire_1208), .Cout(wire_1209),  .A(wire_749), .B(wire_808), .Cin(wire_807));
wire wire_1210, wire_1211;
bit_adder add559(.S(wire_1210), .Cout(wire_1211),  .A(wire_751), .B(wire_810), .Cin(wire_809));
wire wire_1212, wire_1213;
bit_adder add560(.S(wire_1212), .Cout(wire_1213),  .A(wire_753), .B(wire_812), .Cin(wire_811));
wire wire_1214, wire_1215;
bit_adder add561(.S(wire_1214), .Cout(wire_1215),  .A(wire_755), .B(wire_814), .Cin(wire_813));
wire wire_1216, wire_1217;
bit_adder add562(.S(wire_1216), .Cout(wire_1217),  .A(wire_757), .B(wire_816), .Cin(wire_815));
wire wire_1218, wire_1219;
bit_adder add563(.S(wire_1218), .Cout(wire_1219),  .A(wire_759), .B(wire_818), .Cin(wire_817));
wire wire_1220, wire_1221;
bit_adder add564(.S(wire_1220), .Cout(wire_1221),  .A(wire_761), .B(wire_820), .Cin(wire_819));
wire wire_1222, wire_1223;
bit_adder add565(.S(wire_1222), .Cout(wire_1223),  .A(wire_763), .B(wire_822), .Cin(wire_821));
wire wire_1224, wire_1225;
bit_adder add566(.S(wire_1224), .Cout(wire_1225),  .A(wire_765), .B(wire_824), .Cin(wire_823));
wire wire_1226, wire_1227;
bit_adder add567(.S(wire_1226), .Cout(wire_1227),  .A(wire_767), .B(wire_826), .Cin(wire_825));
wire wire_1228, wire_1229;
bit_adder add568(.S(wire_1228), .Cout(wire_1229),  .A(wire_769), .B(wire_828), .Cin(wire_827));
wire wire_1230, wire_1231;
bit_adder add569(.S(wire_1230), .Cout(wire_1231),  .A(wire_771), .B(wire_830), .Cin(wire_829));
wire wire_1232, wire_1233;
assign wire_1232 = wire_832 ^ wire_831;
assign wire_1233 = wire_832 & wire_831;
wire wire_1234, wire_1235;
assign wire_1234 = wire_834 ^ wire_833;
assign wire_1235 = wire_834 & wire_833;
wire wire_1236, wire_1237;
assign wire_1236 = wire_316 ^ wire_835;
assign wire_1237 = wire_316 & wire_835;
wire wire_1238, wire_1239;
assign wire_1238 = wire_838 ^ wire_837;
assign wire_1239 = wire_838 & wire_837;
wire wire_1240, wire_1241;
assign wire_1240 = wire_840 ^ wire_839;
assign wire_1241 = wire_840 & wire_839;
wire wire_1242, wire_1243;
bit_adder add570(.S(wire_1242), .Cout(wire_1243),  .A(wire_842), .B(wire_841), .Cin(partialProduct_18[0]));
wire wire_1244, wire_1245;
bit_adder add571(.S(wire_1244), .Cout(wire_1245),  .A(wire_844), .B(wire_843), .Cin(wire_384));
wire wire_1246, wire_1247;
bit_adder add572(.S(wire_1246), .Cout(wire_1247),  .A(wire_846), .B(wire_845), .Cin(wire_904));
wire wire_1248, wire_1249;
bit_adder add573(.S(wire_1248), .Cout(wire_1249),  .A(wire_848), .B(wire_847), .Cin(wire_906));
wire wire_1250, wire_1251;
bit_adder add574(.S(wire_1250), .Cout(wire_1251),  .A(wire_850), .B(wire_849), .Cin(wire_908));
wire wire_1252, wire_1253;
bit_adder add575(.S(wire_1252), .Cout(wire_1253),  .A(wire_852), .B(wire_851), .Cin(wire_910));
wire wire_1254, wire_1255;
bit_adder add576(.S(wire_1254), .Cout(wire_1255),  .A(wire_854), .B(wire_853), .Cin(wire_912));
wire wire_1256, wire_1257;
bit_adder add577(.S(wire_1256), .Cout(wire_1257),  .A(wire_856), .B(wire_855), .Cin(wire_914));
wire wire_1258, wire_1259;
bit_adder add578(.S(wire_1258), .Cout(wire_1259),  .A(wire_858), .B(wire_857), .Cin(wire_916));
wire wire_1260, wire_1261;
bit_adder add579(.S(wire_1260), .Cout(wire_1261),  .A(wire_860), .B(wire_859), .Cin(wire_918));
wire wire_1262, wire_1263;
bit_adder add580(.S(wire_1262), .Cout(wire_1263),  .A(wire_862), .B(wire_861), .Cin(wire_920));
wire wire_1264, wire_1265;
bit_adder add581(.S(wire_1264), .Cout(wire_1265),  .A(wire_864), .B(wire_863), .Cin(wire_922));
wire wire_1266, wire_1267;
bit_adder add582(.S(wire_1266), .Cout(wire_1267),  .A(wire_866), .B(wire_865), .Cin(wire_924));
wire wire_1268, wire_1269;
bit_adder add583(.S(wire_1268), .Cout(wire_1269),  .A(wire_868), .B(wire_867), .Cin(wire_926));
wire wire_1270, wire_1271;
bit_adder add584(.S(wire_1270), .Cout(wire_1271),  .A(wire_870), .B(wire_869), .Cin(wire_928));
wire wire_1272, wire_1273;
bit_adder add585(.S(wire_1272), .Cout(wire_1273),  .A(wire_872), .B(wire_871), .Cin(wire_930));
wire wire_1274, wire_1275;
bit_adder add586(.S(wire_1274), .Cout(wire_1275),  .A(wire_874), .B(wire_873), .Cin(wire_932));
wire wire_1276, wire_1277;
bit_adder add587(.S(wire_1276), .Cout(wire_1277),  .A(wire_876), .B(wire_875), .Cin(wire_934));
wire wire_1278, wire_1279;
bit_adder add588(.S(wire_1278), .Cout(wire_1279),  .A(wire_878), .B(wire_877), .Cin(wire_936));
wire wire_1280, wire_1281;
bit_adder add589(.S(wire_1280), .Cout(wire_1281),  .A(wire_880), .B(wire_879), .Cin(wire_938));
wire wire_1282, wire_1283;
bit_adder add590(.S(wire_1282), .Cout(wire_1283),  .A(wire_882), .B(wire_881), .Cin(wire_940));
wire wire_1284, wire_1285;
bit_adder add591(.S(wire_1284), .Cout(wire_1285),  .A(wire_884), .B(wire_883), .Cin(wire_942));
wire wire_1286, wire_1287;
bit_adder add592(.S(wire_1286), .Cout(wire_1287),  .A(wire_886), .B(wire_885), .Cin(wire_944));
wire wire_1288, wire_1289;
bit_adder add593(.S(wire_1288), .Cout(wire_1289),  .A(wire_888), .B(wire_887), .Cin(wire_946));
wire wire_1290, wire_1291;
bit_adder add594(.S(wire_1290), .Cout(wire_1291),  .A(wire_890), .B(wire_889), .Cin(wire_948));
wire wire_1292, wire_1293;
bit_adder add595(.S(wire_1292), .Cout(wire_1293),  .A(wire_892), .B(wire_891), .Cin(wire_950));
wire wire_1294, wire_1295;
bit_adder add596(.S(wire_1294), .Cout(wire_1295),  .A(wire_894), .B(wire_893), .Cin(wire_952));
wire wire_1296, wire_1297;
bit_adder add597(.S(wire_1296), .Cout(wire_1297),  .A(wire_896), .B(wire_895), .Cin(wire_954));
wire wire_1298, wire_1299;
bit_adder add598(.S(wire_1298), .Cout(wire_1299),  .A(wire_898), .B(wire_897), .Cin(wire_956));
wire wire_1300, wire_1301;
bit_adder add599(.S(wire_1300), .Cout(wire_1301),  .A(wire_900), .B(wire_899), .Cin(wire_958));
wire wire_1302, wire_1303;
bit_adder add600(.S(wire_1302), .Cout(wire_1303),  .A(wire_902), .B(wire_901), .Cin(wire_960));
wire wire_1304, wire_1305;
assign wire_1304 = wire_903 ^ wire_962;
assign wire_1305 = wire_903 & wire_962;
wire wire_1306, wire_1307;
assign wire_1306 = wire_909 ^ wire_449;
assign wire_1307 = wire_909 & wire_449;
wire wire_1308, wire_1309;
assign wire_1308 = wire_911 ^ wire_968;
assign wire_1309 = wire_911 & wire_968;
wire wire_1310, wire_1311;
bit_adder add601(.S(wire_1310), .Cout(wire_1311),  .A(wire_913), .B(wire_970), .Cin(wire_969));
wire wire_1312, wire_1313;
bit_adder add602(.S(wire_1312), .Cout(wire_1313),  .A(wire_915), .B(wire_972), .Cin(wire_971));
wire wire_1314, wire_1315;
bit_adder add603(.S(wire_1314), .Cout(wire_1315),  .A(wire_917), .B(wire_974), .Cin(wire_973));
wire wire_1316, wire_1317;
bit_adder add604(.S(wire_1316), .Cout(wire_1317),  .A(wire_919), .B(wire_976), .Cin(wire_975));
wire wire_1318, wire_1319;
bit_adder add605(.S(wire_1318), .Cout(wire_1319),  .A(wire_921), .B(wire_978), .Cin(wire_977));
wire wire_1320, wire_1321;
bit_adder add606(.S(wire_1320), .Cout(wire_1321),  .A(wire_923), .B(wire_980), .Cin(wire_979));
wire wire_1322, wire_1323;
bit_adder add607(.S(wire_1322), .Cout(wire_1323),  .A(wire_925), .B(wire_982), .Cin(wire_981));
wire wire_1324, wire_1325;
bit_adder add608(.S(wire_1324), .Cout(wire_1325),  .A(wire_927), .B(wire_984), .Cin(wire_983));
wire wire_1326, wire_1327;
bit_adder add609(.S(wire_1326), .Cout(wire_1327),  .A(wire_929), .B(wire_986), .Cin(wire_985));
wire wire_1328, wire_1329;
bit_adder add610(.S(wire_1328), .Cout(wire_1329),  .A(wire_931), .B(wire_988), .Cin(wire_987));
wire wire_1330, wire_1331;
bit_adder add611(.S(wire_1330), .Cout(wire_1331),  .A(wire_933), .B(wire_990), .Cin(wire_989));
wire wire_1332, wire_1333;
bit_adder add612(.S(wire_1332), .Cout(wire_1333),  .A(wire_935), .B(wire_992), .Cin(wire_991));
wire wire_1334, wire_1335;
bit_adder add613(.S(wire_1334), .Cout(wire_1335),  .A(wire_937), .B(wire_994), .Cin(wire_993));
wire wire_1336, wire_1337;
bit_adder add614(.S(wire_1336), .Cout(wire_1337),  .A(wire_939), .B(wire_996), .Cin(wire_995));
wire wire_1338, wire_1339;
bit_adder add615(.S(wire_1338), .Cout(wire_1339),  .A(wire_941), .B(wire_998), .Cin(wire_997));
wire wire_1340, wire_1341;
bit_adder add616(.S(wire_1340), .Cout(wire_1341),  .A(wire_943), .B(wire_1000), .Cin(wire_999));
wire wire_1342, wire_1343;
bit_adder add617(.S(wire_1342), .Cout(wire_1343),  .A(wire_945), .B(wire_1002), .Cin(wire_1001));
wire wire_1344, wire_1345;
bit_adder add618(.S(wire_1344), .Cout(wire_1345),  .A(wire_947), .B(wire_1004), .Cin(wire_1003));
wire wire_1346, wire_1347;
bit_adder add619(.S(wire_1346), .Cout(wire_1347),  .A(wire_949), .B(wire_1006), .Cin(wire_1005));
wire wire_1348, wire_1349;
bit_adder add620(.S(wire_1348), .Cout(wire_1349),  .A(wire_951), .B(wire_1008), .Cin(wire_1007));
wire wire_1350, wire_1351;
bit_adder add621(.S(wire_1350), .Cout(wire_1351),  .A(wire_953), .B(wire_1010), .Cin(wire_1009));
wire wire_1352, wire_1353;
bit_adder add622(.S(wire_1352), .Cout(wire_1353),  .A(wire_955), .B(wire_1012), .Cin(wire_1011));
wire wire_1354, wire_1355;
bit_adder add623(.S(wire_1354), .Cout(wire_1355),  .A(wire_957), .B(wire_1014), .Cin(wire_1013));
wire wire_1356, wire_1357;
bit_adder add624(.S(wire_1356), .Cout(wire_1357),  .A(wire_959), .B(wire_1016), .Cin(wire_1015));
wire wire_1358, wire_1359;
bit_adder add625(.S(wire_1358), .Cout(wire_1359),  .A(wire_961), .B(wire_1018), .Cin(wire_1017));
wire wire_1360, wire_1361;
bit_adder add626(.S(wire_1360), .Cout(wire_1361),  .A(wire_963), .B(wire_1020), .Cin(wire_1019));
wire wire_1362, wire_1363;
bit_adder add627(.S(wire_1362), .Cout(wire_1363),  .A(wire_965), .B(wire_1022), .Cin(wire_1021));
wire wire_1364, wire_1365;
bit_adder add628(.S(wire_1364), .Cout(wire_1365),  .A(wire_967), .B(wire_1024), .Cin(wire_1023));
wire wire_1366, wire_1367;
assign wire_1366 = wire_1026 ^ wire_1025;
assign wire_1367 = wire_1026 & wire_1025;
wire wire_1368, wire_1369;
assign wire_1368 = wire_1028 ^ wire_1027;
assign wire_1369 = wire_1028 & wire_1027;
wire wire_1370, wire_1371;
assign wire_1370 = wire_1030 ^ wire_1029;
assign wire_1371 = wire_1030 & wire_1029;
wire wire_1372, wire_1373;
assign wire_1372 = wire_1032 ^ wire_1031;
assign wire_1373 = wire_1032 & wire_1031;
wire wire_1374, wire_1375;
assign wire_1374 = wire_1034 ^ wire_1033;
assign wire_1375 = wire_1034 & wire_1033;
wire wire_1376, wire_1377;
assign wire_1376 = wire_1038 ^ wire_1037;
assign wire_1377 = wire_1038 & wire_1037;
wire wire_1378, wire_1379;
bit_adder add629(.S(wire_1378), .Cout(wire_1379),  .A(wire_1040), .B(wire_1039), .Cin(partialProduct_31[0]));
wire wire_1380, wire_1381;
bit_adder add630(.S(wire_1380), .Cout(wire_1381),  .A(wire_1042), .B(wire_1041), .Cin(partialProduct_31[1]));
wire wire_1382, wire_1383;
bit_adder add631(.S(wire_1382), .Cout(wire_1383),  .A(wire_1044), .B(wire_1043), .Cin(partialProduct_31[2]));
wire wire_1384, wire_1385;
bit_adder add632(.S(wire_1384), .Cout(wire_1385),  .A(wire_1046), .B(wire_1045), .Cin(partialProduct_31[3]));
wire wire_1386, wire_1387;
bit_adder add633(.S(wire_1386), .Cout(wire_1387),  .A(wire_1048), .B(wire_1047), .Cin(partialProduct_31[4]));
wire wire_1388, wire_1389;
bit_adder add634(.S(wire_1388), .Cout(wire_1389),  .A(wire_1050), .B(wire_1049), .Cin(partialProduct_31[5]));
wire wire_1390, wire_1391;
bit_adder add635(.S(wire_1390), .Cout(wire_1391),  .A(wire_1052), .B(wire_1051), .Cin(partialProduct_31[6]));
wire wire_1392, wire_1393;
bit_adder add636(.S(wire_1392), .Cout(wire_1393),  .A(wire_1054), .B(wire_1053), .Cin(partialProduct_31[7]));
wire wire_1394, wire_1395;
bit_adder add637(.S(wire_1394), .Cout(wire_1395),  .A(wire_1056), .B(wire_1055), .Cin(partialProduct_31[8]));
wire wire_1396, wire_1397;
bit_adder add638(.S(wire_1396), .Cout(wire_1397),  .A(wire_1058), .B(wire_1057), .Cin(partialProduct_31[9]));
wire wire_1398, wire_1399;
bit_adder add639(.S(wire_1398), .Cout(wire_1399),  .A(wire_1060), .B(wire_1059), .Cin(partialProduct_31[10]));
wire wire_1400, wire_1401;
bit_adder add640(.S(wire_1400), .Cout(wire_1401),  .A(wire_1062), .B(wire_1061), .Cin(partialProduct_31[11]));
wire wire_1402, wire_1403;
bit_adder add641(.S(wire_1402), .Cout(wire_1403),  .A(wire_1064), .B(wire_1063), .Cin(partialProduct_31[12]));
wire wire_1404, wire_1405;
bit_adder add642(.S(wire_1404), .Cout(wire_1405),  .A(wire_1066), .B(wire_1065), .Cin(partialProduct_31[13]));
wire wire_1406, wire_1407;
bit_adder add643(.S(wire_1406), .Cout(wire_1407),  .A(wire_1068), .B(wire_1067), .Cin(partialProduct_31[14]));
wire wire_1408, wire_1409;
bit_adder add644(.S(wire_1408), .Cout(wire_1409),  .A(wire_1070), .B(wire_1069), .Cin(partialProduct_31[15]));
wire wire_1410, wire_1411;
bit_adder add645(.S(wire_1410), .Cout(wire_1411),  .A(wire_1072), .B(wire_1071), .Cin(partialProduct_31[16]));
wire wire_1412, wire_1413;
bit_adder add646(.S(wire_1412), .Cout(wire_1413),  .A(wire_1074), .B(wire_1073), .Cin(partialProduct_31[17]));
wire wire_1414, wire_1415;
bit_adder add647(.S(wire_1414), .Cout(wire_1415),  .A(wire_1076), .B(wire_1075), .Cin(partialProduct_31[18]));
wire wire_1416, wire_1417;
bit_adder add648(.S(wire_1416), .Cout(wire_1417),  .A(wire_1078), .B(wire_1077), .Cin(partialProduct_31[19]));
wire wire_1418, wire_1419;
bit_adder add649(.S(wire_1418), .Cout(wire_1419),  .A(wire_1080), .B(wire_1079), .Cin(partialProduct_31[20]));
wire wire_1420, wire_1421;
bit_adder add650(.S(wire_1420), .Cout(wire_1421),  .A(wire_1082), .B(wire_1081), .Cin(partialProduct_31[21]));
wire wire_1422, wire_1423;
bit_adder add651(.S(wire_1422), .Cout(wire_1423),  .A(wire_1084), .B(wire_1083), .Cin(partialProduct_31[22]));
wire wire_1424, wire_1425;
bit_adder add652(.S(wire_1424), .Cout(wire_1425),  .A(wire_1086), .B(wire_1085), .Cin(partialProduct_31[23]));
wire wire_1426, wire_1427;
bit_adder add653(.S(wire_1426), .Cout(wire_1427),  .A(wire_1088), .B(wire_1087), .Cin(partialProduct_31[24]));
wire wire_1428, wire_1429;
bit_adder add654(.S(wire_1428), .Cout(wire_1429),  .A(wire_1090), .B(wire_1089), .Cin(partialProduct_31[25]));
wire wire_1430, wire_1431;
bit_adder add655(.S(wire_1430), .Cout(wire_1431),  .A(wire_1092), .B(wire_1091), .Cin(partialProduct_31[26]));
wire wire_1432, wire_1433;
bit_adder add656(.S(wire_1432), .Cout(wire_1433),  .A(wire_1094), .B(wire_1093), .Cin(partialProduct_31[27]));
wire wire_1434, wire_1435;
bit_adder add657(.S(wire_1434), .Cout(wire_1435),  .A(wire_1096), .B(wire_1095), .Cin(partialProduct_31[28]));
wire wire_1436, wire_1437;
bit_adder add658(.S(wire_1436), .Cout(wire_1437),  .A(wire_1098), .B(wire_1097), .Cin(partialProduct_31[29]));
wire wire_1438, wire_1439;
bit_adder add659(.S(wire_1438), .Cout(wire_1439),  .A(partialProduct_30[31]), .B(wire_1099), .Cin(partialProduct_31[30]));
wire wire_1440, wire_1441;
assign wire_1440 = wire_1102 ^ wire_1101;
assign wire_1441 = wire_1102 & wire_1101;
wire wire_1442, wire_1443;
assign wire_1442 = wire_1104 ^ wire_1103;
assign wire_1443 = wire_1104 & wire_1103;
wire wire_1444, wire_1445;
assign wire_1444 = wire_1106 ^ wire_1105;
assign wire_1445 = wire_1106 & wire_1105;
wire wire_1446, wire_1447;
bit_adder add660(.S(wire_1446), .Cout(wire_1447),  .A(wire_1108), .B(wire_1107), .Cin(wire_705));
wire wire_1448, wire_1449;
bit_adder add661(.S(wire_1448), .Cout(wire_1449),  .A(wire_1110), .B(wire_1109), .Cin(wire_707));
wire wire_1450, wire_1451;
bit_adder add662(.S(wire_1450), .Cout(wire_1451),  .A(wire_1112), .B(wire_1111), .Cin(wire_1168));
wire wire_1452, wire_1453;
bit_adder add663(.S(wire_1452), .Cout(wire_1453),  .A(wire_1114), .B(wire_1113), .Cin(wire_1170));
wire wire_1454, wire_1455;
bit_adder add664(.S(wire_1454), .Cout(wire_1455),  .A(wire_1116), .B(wire_1115), .Cin(wire_1172));
wire wire_1456, wire_1457;
bit_adder add665(.S(wire_1456), .Cout(wire_1457),  .A(wire_1118), .B(wire_1117), .Cin(wire_1174));
wire wire_1458, wire_1459;
bit_adder add666(.S(wire_1458), .Cout(wire_1459),  .A(wire_1120), .B(wire_1119), .Cin(wire_1176));
wire wire_1460, wire_1461;
bit_adder add667(.S(wire_1460), .Cout(wire_1461),  .A(wire_1122), .B(wire_1121), .Cin(wire_1178));
wire wire_1462, wire_1463;
bit_adder add668(.S(wire_1462), .Cout(wire_1463),  .A(wire_1124), .B(wire_1123), .Cin(wire_1180));
wire wire_1464, wire_1465;
bit_adder add669(.S(wire_1464), .Cout(wire_1465),  .A(wire_1126), .B(wire_1125), .Cin(wire_1182));
wire wire_1466, wire_1467;
bit_adder add670(.S(wire_1466), .Cout(wire_1467),  .A(wire_1128), .B(wire_1127), .Cin(wire_1184));
wire wire_1468, wire_1469;
bit_adder add671(.S(wire_1468), .Cout(wire_1469),  .A(wire_1130), .B(wire_1129), .Cin(wire_1186));
wire wire_1470, wire_1471;
bit_adder add672(.S(wire_1470), .Cout(wire_1471),  .A(wire_1132), .B(wire_1131), .Cin(wire_1188));
wire wire_1472, wire_1473;
bit_adder add673(.S(wire_1472), .Cout(wire_1473),  .A(wire_1134), .B(wire_1133), .Cin(wire_1190));
wire wire_1474, wire_1475;
bit_adder add674(.S(wire_1474), .Cout(wire_1475),  .A(wire_1136), .B(wire_1135), .Cin(wire_1192));
wire wire_1476, wire_1477;
bit_adder add675(.S(wire_1476), .Cout(wire_1477),  .A(wire_1138), .B(wire_1137), .Cin(wire_1194));
wire wire_1478, wire_1479;
bit_adder add676(.S(wire_1478), .Cout(wire_1479),  .A(wire_1140), .B(wire_1139), .Cin(wire_1196));
wire wire_1480, wire_1481;
bit_adder add677(.S(wire_1480), .Cout(wire_1481),  .A(wire_1142), .B(wire_1141), .Cin(wire_1198));
wire wire_1482, wire_1483;
bit_adder add678(.S(wire_1482), .Cout(wire_1483),  .A(wire_1144), .B(wire_1143), .Cin(wire_1200));
wire wire_1484, wire_1485;
bit_adder add679(.S(wire_1484), .Cout(wire_1485),  .A(wire_1146), .B(wire_1145), .Cin(wire_1202));
wire wire_1486, wire_1487;
bit_adder add680(.S(wire_1486), .Cout(wire_1487),  .A(wire_1148), .B(wire_1147), .Cin(wire_1204));
wire wire_1488, wire_1489;
bit_adder add681(.S(wire_1488), .Cout(wire_1489),  .A(wire_1150), .B(wire_1149), .Cin(wire_1206));
wire wire_1490, wire_1491;
bit_adder add682(.S(wire_1490), .Cout(wire_1491),  .A(wire_1152), .B(wire_1151), .Cin(wire_1208));
wire wire_1492, wire_1493;
bit_adder add683(.S(wire_1492), .Cout(wire_1493),  .A(wire_1154), .B(wire_1153), .Cin(wire_1210));
wire wire_1494, wire_1495;
bit_adder add684(.S(wire_1494), .Cout(wire_1495),  .A(wire_1156), .B(wire_1155), .Cin(wire_1212));
wire wire_1496, wire_1497;
bit_adder add685(.S(wire_1496), .Cout(wire_1497),  .A(wire_1158), .B(wire_1157), .Cin(wire_1214));
wire wire_1498, wire_1499;
bit_adder add686(.S(wire_1498), .Cout(wire_1499),  .A(wire_1160), .B(wire_1159), .Cin(wire_1216));
wire wire_1500, wire_1501;
bit_adder add687(.S(wire_1500), .Cout(wire_1501),  .A(wire_1162), .B(wire_1161), .Cin(wire_1218));
wire wire_1502, wire_1503;
bit_adder add688(.S(wire_1502), .Cout(wire_1503),  .A(wire_1164), .B(wire_1163), .Cin(wire_1220));
wire wire_1504, wire_1505;
bit_adder add689(.S(wire_1504), .Cout(wire_1505),  .A(wire_1166), .B(wire_1165), .Cin(wire_1222));
wire wire_1506, wire_1507;
bit_adder add690(.S(wire_1506), .Cout(wire_1507),  .A(wire_766), .B(wire_1167), .Cin(wire_1224));
wire wire_1508, wire_1509;
assign wire_1508 = wire_768 ^ wire_1226;
assign wire_1509 = wire_768 & wire_1226;
wire wire_1510, wire_1511;
assign wire_1510 = wire_770 ^ wire_1228;
assign wire_1511 = wire_770 & wire_1228;
wire wire_1512, wire_1513;
assign wire_1512 = wire_1177 ^ wire_257;
assign wire_1513 = wire_1177 & wire_257;
wire wire_1514, wire_1515;
assign wire_1514 = wire_1179 ^ wire_836;
assign wire_1515 = wire_1179 & wire_836;
wire wire_1516, wire_1517;
assign wire_1516 = wire_1181 ^ wire_1238;
assign wire_1517 = wire_1181 & wire_1238;
wire wire_1518, wire_1519;
bit_adder add691(.S(wire_1518), .Cout(wire_1519),  .A(wire_1183), .B(wire_1240), .Cin(wire_1239));
wire wire_1520, wire_1521;
bit_adder add692(.S(wire_1520), .Cout(wire_1521),  .A(wire_1185), .B(wire_1242), .Cin(wire_1241));
wire wire_1522, wire_1523;
bit_adder add693(.S(wire_1522), .Cout(wire_1523),  .A(wire_1187), .B(wire_1244), .Cin(wire_1243));
wire wire_1524, wire_1525;
bit_adder add694(.S(wire_1524), .Cout(wire_1525),  .A(wire_1189), .B(wire_1246), .Cin(wire_1245));
wire wire_1526, wire_1527;
bit_adder add695(.S(wire_1526), .Cout(wire_1527),  .A(wire_1191), .B(wire_1248), .Cin(wire_1247));
wire wire_1528, wire_1529;
bit_adder add696(.S(wire_1528), .Cout(wire_1529),  .A(wire_1193), .B(wire_1250), .Cin(wire_1249));
wire wire_1530, wire_1531;
bit_adder add697(.S(wire_1530), .Cout(wire_1531),  .A(wire_1195), .B(wire_1252), .Cin(wire_1251));
wire wire_1532, wire_1533;
bit_adder add698(.S(wire_1532), .Cout(wire_1533),  .A(wire_1197), .B(wire_1254), .Cin(wire_1253));
wire wire_1534, wire_1535;
bit_adder add699(.S(wire_1534), .Cout(wire_1535),  .A(wire_1199), .B(wire_1256), .Cin(wire_1255));
wire wire_1536, wire_1537;
bit_adder add700(.S(wire_1536), .Cout(wire_1537),  .A(wire_1201), .B(wire_1258), .Cin(wire_1257));
wire wire_1538, wire_1539;
bit_adder add701(.S(wire_1538), .Cout(wire_1539),  .A(wire_1203), .B(wire_1260), .Cin(wire_1259));
wire wire_1540, wire_1541;
bit_adder add702(.S(wire_1540), .Cout(wire_1541),  .A(wire_1205), .B(wire_1262), .Cin(wire_1261));
wire wire_1542, wire_1543;
bit_adder add703(.S(wire_1542), .Cout(wire_1543),  .A(wire_1207), .B(wire_1264), .Cin(wire_1263));
wire wire_1544, wire_1545;
bit_adder add704(.S(wire_1544), .Cout(wire_1545),  .A(wire_1209), .B(wire_1266), .Cin(wire_1265));
wire wire_1546, wire_1547;
bit_adder add705(.S(wire_1546), .Cout(wire_1547),  .A(wire_1211), .B(wire_1268), .Cin(wire_1267));
wire wire_1548, wire_1549;
bit_adder add706(.S(wire_1548), .Cout(wire_1549),  .A(wire_1213), .B(wire_1270), .Cin(wire_1269));
wire wire_1550, wire_1551;
bit_adder add707(.S(wire_1550), .Cout(wire_1551),  .A(wire_1215), .B(wire_1272), .Cin(wire_1271));
wire wire_1552, wire_1553;
bit_adder add708(.S(wire_1552), .Cout(wire_1553),  .A(wire_1217), .B(wire_1274), .Cin(wire_1273));
wire wire_1554, wire_1555;
bit_adder add709(.S(wire_1554), .Cout(wire_1555),  .A(wire_1219), .B(wire_1276), .Cin(wire_1275));
wire wire_1556, wire_1557;
bit_adder add710(.S(wire_1556), .Cout(wire_1557),  .A(wire_1221), .B(wire_1278), .Cin(wire_1277));
wire wire_1558, wire_1559;
bit_adder add711(.S(wire_1558), .Cout(wire_1559),  .A(wire_1223), .B(wire_1280), .Cin(wire_1279));
wire wire_1560, wire_1561;
bit_adder add712(.S(wire_1560), .Cout(wire_1561),  .A(wire_1225), .B(wire_1282), .Cin(wire_1281));
wire wire_1562, wire_1563;
bit_adder add713(.S(wire_1562), .Cout(wire_1563),  .A(wire_1227), .B(wire_1284), .Cin(wire_1283));
wire wire_1564, wire_1565;
bit_adder add714(.S(wire_1564), .Cout(wire_1565),  .A(wire_1229), .B(wire_1286), .Cin(wire_1285));
wire wire_1566, wire_1567;
bit_adder add715(.S(wire_1566), .Cout(wire_1567),  .A(wire_1231), .B(wire_1288), .Cin(wire_1287));
wire wire_1568, wire_1569;
bit_adder add716(.S(wire_1568), .Cout(wire_1569),  .A(wire_1233), .B(wire_1290), .Cin(wire_1289));
wire wire_1570, wire_1571;
bit_adder add717(.S(wire_1570), .Cout(wire_1571),  .A(wire_1235), .B(wire_1292), .Cin(wire_1291));
wire wire_1572, wire_1573;
bit_adder add718(.S(wire_1572), .Cout(wire_1573),  .A(wire_1237), .B(wire_1294), .Cin(wire_1293));
wire wire_1574, wire_1575;
assign wire_1574 = wire_1296 ^ wire_1295;
assign wire_1575 = wire_1296 & wire_1295;
wire wire_1576, wire_1577;
assign wire_1576 = wire_1298 ^ wire_1297;
assign wire_1577 = wire_1298 & wire_1297;
wire wire_1578, wire_1579;
assign wire_1578 = wire_1300 ^ wire_1299;
assign wire_1579 = wire_1300 & wire_1299;
wire wire_1580, wire_1581;
assign wire_1580 = wire_1302 ^ wire_1301;
assign wire_1581 = wire_1302 & wire_1301;
wire wire_1582, wire_1583;
assign wire_1582 = wire_1304 ^ wire_1303;
assign wire_1583 = wire_1304 & wire_1303;
wire wire_1584, wire_1585;
assign wire_1584 = wire_964 ^ wire_1305;
assign wire_1585 = wire_964 & wire_1305;
wire wire_1586, wire_1587;
assign wire_1586 = wire_1308 ^ wire_1307;
assign wire_1587 = wire_1308 & wire_1307;
wire wire_1588, wire_1589;
assign wire_1588 = wire_1310 ^ wire_1309;
assign wire_1589 = wire_1310 & wire_1309;
wire wire_1590, wire_1591;
assign wire_1590 = wire_1312 ^ wire_1311;
assign wire_1591 = wire_1312 & wire_1311;
wire wire_1592, wire_1593;
bit_adder add719(.S(wire_1592), .Cout(wire_1593),  .A(wire_1314), .B(wire_1313), .Cin(partialProduct_27[0]));
wire wire_1594, wire_1595;
bit_adder add720(.S(wire_1594), .Cout(wire_1595),  .A(wire_1316), .B(wire_1315), .Cin(wire_576));
wire wire_1596, wire_1597;
bit_adder add721(.S(wire_1596), .Cout(wire_1597),  .A(wire_1318), .B(wire_1317), .Cin(wire_1036));
wire wire_1598, wire_1599;
bit_adder add722(.S(wire_1598), .Cout(wire_1599),  .A(wire_1320), .B(wire_1319), .Cin(wire_1376));
wire wire_1600, wire_1601;
bit_adder add723(.S(wire_1600), .Cout(wire_1601),  .A(wire_1322), .B(wire_1321), .Cin(wire_1378));
wire wire_1602, wire_1603;
bit_adder add724(.S(wire_1602), .Cout(wire_1603),  .A(wire_1324), .B(wire_1323), .Cin(wire_1380));
wire wire_1604, wire_1605;
bit_adder add725(.S(wire_1604), .Cout(wire_1605),  .A(wire_1326), .B(wire_1325), .Cin(wire_1382));
wire wire_1606, wire_1607;
bit_adder add726(.S(wire_1606), .Cout(wire_1607),  .A(wire_1328), .B(wire_1327), .Cin(wire_1384));
wire wire_1608, wire_1609;
bit_adder add727(.S(wire_1608), .Cout(wire_1609),  .A(wire_1330), .B(wire_1329), .Cin(wire_1386));
wire wire_1610, wire_1611;
bit_adder add728(.S(wire_1610), .Cout(wire_1611),  .A(wire_1332), .B(wire_1331), .Cin(wire_1388));
wire wire_1612, wire_1613;
bit_adder add729(.S(wire_1612), .Cout(wire_1613),  .A(wire_1334), .B(wire_1333), .Cin(wire_1390));
wire wire_1614, wire_1615;
bit_adder add730(.S(wire_1614), .Cout(wire_1615),  .A(wire_1336), .B(wire_1335), .Cin(wire_1392));
wire wire_1616, wire_1617;
bit_adder add731(.S(wire_1616), .Cout(wire_1617),  .A(wire_1338), .B(wire_1337), .Cin(wire_1394));
wire wire_1618, wire_1619;
bit_adder add732(.S(wire_1618), .Cout(wire_1619),  .A(wire_1340), .B(wire_1339), .Cin(wire_1396));
wire wire_1620, wire_1621;
bit_adder add733(.S(wire_1620), .Cout(wire_1621),  .A(wire_1342), .B(wire_1341), .Cin(wire_1398));
wire wire_1622, wire_1623;
bit_adder add734(.S(wire_1622), .Cout(wire_1623),  .A(wire_1344), .B(wire_1343), .Cin(wire_1400));
wire wire_1624, wire_1625;
bit_adder add735(.S(wire_1624), .Cout(wire_1625),  .A(wire_1346), .B(wire_1345), .Cin(wire_1402));
wire wire_1626, wire_1627;
bit_adder add736(.S(wire_1626), .Cout(wire_1627),  .A(wire_1348), .B(wire_1347), .Cin(wire_1404));
wire wire_1628, wire_1629;
bit_adder add737(.S(wire_1628), .Cout(wire_1629),  .A(wire_1350), .B(wire_1349), .Cin(wire_1406));
wire wire_1630, wire_1631;
bit_adder add738(.S(wire_1630), .Cout(wire_1631),  .A(wire_1352), .B(wire_1351), .Cin(wire_1408));
wire wire_1632, wire_1633;
bit_adder add739(.S(wire_1632), .Cout(wire_1633),  .A(wire_1354), .B(wire_1353), .Cin(wire_1410));
wire wire_1634, wire_1635;
bit_adder add740(.S(wire_1634), .Cout(wire_1635),  .A(wire_1356), .B(wire_1355), .Cin(wire_1412));
wire wire_1636, wire_1637;
bit_adder add741(.S(wire_1636), .Cout(wire_1637),  .A(wire_1358), .B(wire_1357), .Cin(wire_1414));
wire wire_1638, wire_1639;
bit_adder add742(.S(wire_1638), .Cout(wire_1639),  .A(wire_1360), .B(wire_1359), .Cin(wire_1416));
wire wire_1640, wire_1641;
bit_adder add743(.S(wire_1640), .Cout(wire_1641),  .A(wire_1362), .B(wire_1361), .Cin(wire_1418));
wire wire_1642, wire_1643;
bit_adder add744(.S(wire_1642), .Cout(wire_1643),  .A(wire_1364), .B(wire_1363), .Cin(wire_1420));
wire wire_1644, wire_1645;
bit_adder add745(.S(wire_1644), .Cout(wire_1645),  .A(wire_1366), .B(wire_1365), .Cin(wire_1422));
wire wire_1646, wire_1647;
bit_adder add746(.S(wire_1646), .Cout(wire_1647),  .A(wire_1368), .B(wire_1367), .Cin(wire_1424));
wire wire_1648, wire_1649;
bit_adder add747(.S(wire_1648), .Cout(wire_1649),  .A(wire_1370), .B(wire_1369), .Cin(wire_1426));
wire wire_1650, wire_1651;
bit_adder add748(.S(wire_1650), .Cout(wire_1651),  .A(wire_1372), .B(wire_1371), .Cin(wire_1428));
wire wire_1652, wire_1653;
bit_adder add749(.S(wire_1652), .Cout(wire_1653),  .A(wire_1374), .B(wire_1373), .Cin(wire_1430));
wire wire_1654, wire_1655;
bit_adder add750(.S(wire_1654), .Cout(wire_1655),  .A(wire_1035), .B(wire_1375), .Cin(wire_1432));
wire wire_1656, wire_1657;
assign wire_1656 = wire_1442 ^ wire_1441;
assign wire_1657 = wire_1442 & wire_1441;
wire wire_1658, wire_1659;
assign wire_1658 = wire_1444 ^ wire_1443;
assign wire_1659 = wire_1444 & wire_1443;
wire wire_1660, wire_1661;
assign wire_1660 = wire_1446 ^ wire_1445;
assign wire_1661 = wire_1446 & wire_1445;
wire wire_1662, wire_1663;
assign wire_1662 = wire_1448 ^ wire_1447;
assign wire_1663 = wire_1448 & wire_1447;
wire wire_1664, wire_1665;
assign wire_1664 = wire_1450 ^ wire_1449;
assign wire_1665 = wire_1450 & wire_1449;
wire wire_1666, wire_1667;
bit_adder add751(.S(wire_1666), .Cout(wire_1667),  .A(wire_1452), .B(wire_1451), .Cin(wire_1169));
wire wire_1668, wire_1669;
bit_adder add752(.S(wire_1668), .Cout(wire_1669),  .A(wire_1454), .B(wire_1453), .Cin(wire_1171));
wire wire_1670, wire_1671;
bit_adder add753(.S(wire_1670), .Cout(wire_1671),  .A(wire_1456), .B(wire_1455), .Cin(wire_1173));
wire wire_1672, wire_1673;
bit_adder add754(.S(wire_1672), .Cout(wire_1673),  .A(wire_1458), .B(wire_1457), .Cin(wire_1175));
wire wire_1674, wire_1675;
bit_adder add755(.S(wire_1674), .Cout(wire_1675),  .A(wire_1460), .B(wire_1459), .Cin(wire_1512));
wire wire_1676, wire_1677;
bit_adder add756(.S(wire_1676), .Cout(wire_1677),  .A(wire_1462), .B(wire_1461), .Cin(wire_1514));
wire wire_1678, wire_1679;
bit_adder add757(.S(wire_1678), .Cout(wire_1679),  .A(wire_1464), .B(wire_1463), .Cin(wire_1516));
wire wire_1680, wire_1681;
bit_adder add758(.S(wire_1680), .Cout(wire_1681),  .A(wire_1466), .B(wire_1465), .Cin(wire_1518));
wire wire_1682, wire_1683;
bit_adder add759(.S(wire_1682), .Cout(wire_1683),  .A(wire_1468), .B(wire_1467), .Cin(wire_1520));
wire wire_1684, wire_1685;
bit_adder add760(.S(wire_1684), .Cout(wire_1685),  .A(wire_1470), .B(wire_1469), .Cin(wire_1522));
wire wire_1686, wire_1687;
bit_adder add761(.S(wire_1686), .Cout(wire_1687),  .A(wire_1472), .B(wire_1471), .Cin(wire_1524));
wire wire_1688, wire_1689;
bit_adder add762(.S(wire_1688), .Cout(wire_1689),  .A(wire_1474), .B(wire_1473), .Cin(wire_1526));
wire wire_1690, wire_1691;
bit_adder add763(.S(wire_1690), .Cout(wire_1691),  .A(wire_1476), .B(wire_1475), .Cin(wire_1528));
wire wire_1692, wire_1693;
bit_adder add764(.S(wire_1692), .Cout(wire_1693),  .A(wire_1478), .B(wire_1477), .Cin(wire_1530));
wire wire_1694, wire_1695;
bit_adder add765(.S(wire_1694), .Cout(wire_1695),  .A(wire_1480), .B(wire_1479), .Cin(wire_1532));
wire wire_1696, wire_1697;
bit_adder add766(.S(wire_1696), .Cout(wire_1697),  .A(wire_1482), .B(wire_1481), .Cin(wire_1534));
wire wire_1698, wire_1699;
bit_adder add767(.S(wire_1698), .Cout(wire_1699),  .A(wire_1484), .B(wire_1483), .Cin(wire_1536));
wire wire_1700, wire_1701;
bit_adder add768(.S(wire_1700), .Cout(wire_1701),  .A(wire_1486), .B(wire_1485), .Cin(wire_1538));
wire wire_1702, wire_1703;
bit_adder add769(.S(wire_1702), .Cout(wire_1703),  .A(wire_1488), .B(wire_1487), .Cin(wire_1540));
wire wire_1704, wire_1705;
bit_adder add770(.S(wire_1704), .Cout(wire_1705),  .A(wire_1490), .B(wire_1489), .Cin(wire_1542));
wire wire_1706, wire_1707;
bit_adder add771(.S(wire_1706), .Cout(wire_1707),  .A(wire_1492), .B(wire_1491), .Cin(wire_1544));
wire wire_1708, wire_1709;
bit_adder add772(.S(wire_1708), .Cout(wire_1709),  .A(wire_1494), .B(wire_1493), .Cin(wire_1546));
wire wire_1710, wire_1711;
bit_adder add773(.S(wire_1710), .Cout(wire_1711),  .A(wire_1496), .B(wire_1495), .Cin(wire_1548));
wire wire_1712, wire_1713;
bit_adder add774(.S(wire_1712), .Cout(wire_1713),  .A(wire_1498), .B(wire_1497), .Cin(wire_1550));
wire wire_1714, wire_1715;
bit_adder add775(.S(wire_1714), .Cout(wire_1715),  .A(wire_1500), .B(wire_1499), .Cin(wire_1552));
wire wire_1716, wire_1717;
bit_adder add776(.S(wire_1716), .Cout(wire_1717),  .A(wire_1502), .B(wire_1501), .Cin(wire_1554));
wire wire_1718, wire_1719;
bit_adder add777(.S(wire_1718), .Cout(wire_1719),  .A(wire_1504), .B(wire_1503), .Cin(wire_1556));
wire wire_1720, wire_1721;
bit_adder add778(.S(wire_1720), .Cout(wire_1721),  .A(wire_1506), .B(wire_1505), .Cin(wire_1558));
wire wire_1722, wire_1723;
bit_adder add779(.S(wire_1722), .Cout(wire_1723),  .A(wire_1508), .B(wire_1507), .Cin(wire_1560));
wire wire_1724, wire_1725;
bit_adder add780(.S(wire_1724), .Cout(wire_1725),  .A(wire_1510), .B(wire_1509), .Cin(wire_1562));
wire wire_1726, wire_1727;
bit_adder add781(.S(wire_1726), .Cout(wire_1727),  .A(wire_1230), .B(wire_1511), .Cin(wire_1564));
wire wire_1728, wire_1729;
assign wire_1728 = wire_1232 ^ wire_1566;
assign wire_1729 = wire_1232 & wire_1566;
wire wire_1730, wire_1731;
assign wire_1730 = wire_1234 ^ wire_1568;
assign wire_1731 = wire_1234 & wire_1568;
wire wire_1732, wire_1733;
assign wire_1732 = wire_1236 ^ wire_1570;
assign wire_1733 = wire_1236 & wire_1570;
wire wire_1734, wire_1735;
assign wire_1734 = wire_318 ^ wire_1572;
assign wire_1735 = wire_318 & wire_1572;
wire wire_1736, wire_1737;
assign wire_1736 = partialProduct_14[31] ^ wire_1574;
assign wire_1737 = partialProduct_14[31] & wire_1574;
wire wire_1738, wire_1739;
assign wire_1738 = wire_1525 ^ wire_905;
assign wire_1739 = wire_1525 & wire_905;
wire wire_1740, wire_1741;
assign wire_1740 = wire_1527 ^ wire_907;
assign wire_1741 = wire_1527 & wire_907;
wire wire_1742, wire_1743;
assign wire_1742 = wire_1529 ^ wire_1306;
assign wire_1743 = wire_1529 & wire_1306;
wire wire_1744, wire_1745;
assign wire_1744 = wire_1531 ^ wire_1586;
assign wire_1745 = wire_1531 & wire_1586;
wire wire_1746, wire_1747;
bit_adder add782(.S(wire_1746), .Cout(wire_1747),  .A(wire_1533), .B(wire_1588), .Cin(wire_1587));
wire wire_1748, wire_1749;
bit_adder add783(.S(wire_1748), .Cout(wire_1749),  .A(wire_1535), .B(wire_1590), .Cin(wire_1589));
wire wire_1750, wire_1751;
bit_adder add784(.S(wire_1750), .Cout(wire_1751),  .A(wire_1537), .B(wire_1592), .Cin(wire_1591));
wire wire_1752, wire_1753;
bit_adder add785(.S(wire_1752), .Cout(wire_1753),  .A(wire_1539), .B(wire_1594), .Cin(wire_1593));
wire wire_1754, wire_1755;
bit_adder add786(.S(wire_1754), .Cout(wire_1755),  .A(wire_1541), .B(wire_1596), .Cin(wire_1595));
wire wire_1756, wire_1757;
bit_adder add787(.S(wire_1756), .Cout(wire_1757),  .A(wire_1543), .B(wire_1598), .Cin(wire_1597));
wire wire_1758, wire_1759;
bit_adder add788(.S(wire_1758), .Cout(wire_1759),  .A(wire_1545), .B(wire_1600), .Cin(wire_1599));
wire wire_1760, wire_1761;
bit_adder add789(.S(wire_1760), .Cout(wire_1761),  .A(wire_1547), .B(wire_1602), .Cin(wire_1601));
wire wire_1762, wire_1763;
bit_adder add790(.S(wire_1762), .Cout(wire_1763),  .A(wire_1549), .B(wire_1604), .Cin(wire_1603));
wire wire_1764, wire_1765;
bit_adder add791(.S(wire_1764), .Cout(wire_1765),  .A(wire_1551), .B(wire_1606), .Cin(wire_1605));
wire wire_1766, wire_1767;
bit_adder add792(.S(wire_1766), .Cout(wire_1767),  .A(wire_1553), .B(wire_1608), .Cin(wire_1607));
wire wire_1768, wire_1769;
bit_adder add793(.S(wire_1768), .Cout(wire_1769),  .A(wire_1555), .B(wire_1610), .Cin(wire_1609));
wire wire_1770, wire_1771;
bit_adder add794(.S(wire_1770), .Cout(wire_1771),  .A(wire_1557), .B(wire_1612), .Cin(wire_1611));
wire wire_1772, wire_1773;
bit_adder add795(.S(wire_1772), .Cout(wire_1773),  .A(wire_1559), .B(wire_1614), .Cin(wire_1613));
wire wire_1774, wire_1775;
bit_adder add796(.S(wire_1774), .Cout(wire_1775),  .A(wire_1561), .B(wire_1616), .Cin(wire_1615));
wire wire_1776, wire_1777;
bit_adder add797(.S(wire_1776), .Cout(wire_1777),  .A(wire_1563), .B(wire_1618), .Cin(wire_1617));
wire wire_1778, wire_1779;
bit_adder add798(.S(wire_1778), .Cout(wire_1779),  .A(wire_1565), .B(wire_1620), .Cin(wire_1619));
wire wire_1780, wire_1781;
bit_adder add799(.S(wire_1780), .Cout(wire_1781),  .A(wire_1567), .B(wire_1622), .Cin(wire_1621));
wire wire_1782, wire_1783;
bit_adder add800(.S(wire_1782), .Cout(wire_1783),  .A(wire_1569), .B(wire_1624), .Cin(wire_1623));
wire wire_1784, wire_1785;
bit_adder add801(.S(wire_1784), .Cout(wire_1785),  .A(wire_1571), .B(wire_1626), .Cin(wire_1625));
wire wire_1786, wire_1787;
bit_adder add802(.S(wire_1786), .Cout(wire_1787),  .A(wire_1573), .B(wire_1628), .Cin(wire_1627));
wire wire_1788, wire_1789;
bit_adder add803(.S(wire_1788), .Cout(wire_1789),  .A(wire_1575), .B(wire_1630), .Cin(wire_1629));
wire wire_1790, wire_1791;
bit_adder add804(.S(wire_1790), .Cout(wire_1791),  .A(wire_1577), .B(wire_1632), .Cin(wire_1631));
wire wire_1792, wire_1793;
bit_adder add805(.S(wire_1792), .Cout(wire_1793),  .A(wire_1579), .B(wire_1634), .Cin(wire_1633));
wire wire_1794, wire_1795;
bit_adder add806(.S(wire_1794), .Cout(wire_1795),  .A(wire_1581), .B(wire_1636), .Cin(wire_1635));
wire wire_1796, wire_1797;
bit_adder add807(.S(wire_1796), .Cout(wire_1797),  .A(wire_1583), .B(wire_1638), .Cin(wire_1637));
wire wire_1798, wire_1799;
bit_adder add808(.S(wire_1798), .Cout(wire_1799),  .A(wire_1585), .B(wire_1640), .Cin(wire_1639));
wire wire_1800, wire_1801;
assign wire_1800 = wire_1642 ^ wire_1641;
assign wire_1801 = wire_1642 & wire_1641;
wire wire_1802, wire_1803;
assign wire_1802 = wire_1644 ^ wire_1643;
assign wire_1803 = wire_1644 & wire_1643;
wire wire_1804, wire_1805;
assign wire_1804 = wire_1646 ^ wire_1645;
assign wire_1805 = wire_1646 & wire_1645;
wire wire_1806, wire_1807;
assign wire_1806 = wire_1648 ^ wire_1647;
assign wire_1807 = wire_1648 & wire_1647;
wire wire_1808, wire_1809;
assign wire_1808 = wire_1650 ^ wire_1649;
assign wire_1809 = wire_1650 & wire_1649;
wire wire_1810, wire_1811;
assign wire_1810 = wire_1652 ^ wire_1651;
assign wire_1811 = wire_1652 & wire_1651;
wire wire_1812, wire_1813;
assign wire_1812 = wire_1654 ^ wire_1653;
assign wire_1813 = wire_1654 & wire_1653;
wire wire_1814, wire_1815;
assign wire_1814 = wire_1434 ^ wire_1655;
assign wire_1815 = wire_1434 & wire_1655;
wire wire_1816, wire_1817;
assign wire_1816 = wire_1658 ^ wire_1657;
assign wire_1817 = wire_1658 & wire_1657;
wire wire_1818, wire_1819;
assign wire_1818 = wire_1660 ^ wire_1659;
assign wire_1819 = wire_1660 & wire_1659;
wire wire_1820, wire_1821;
assign wire_1820 = wire_1662 ^ wire_1661;
assign wire_1821 = wire_1662 & wire_1661;
wire wire_1822, wire_1823;
assign wire_1822 = wire_1664 ^ wire_1663;
assign wire_1823 = wire_1664 & wire_1663;
wire wire_1824, wire_1825;
assign wire_1824 = wire_1666 ^ wire_1665;
assign wire_1825 = wire_1666 & wire_1665;
wire wire_1826, wire_1827;
assign wire_1826 = wire_1668 ^ wire_1667;
assign wire_1827 = wire_1668 & wire_1667;
wire wire_1828, wire_1829;
assign wire_1828 = wire_1670 ^ wire_1669;
assign wire_1829 = wire_1670 & wire_1669;
wire wire_1830, wire_1831;
assign wire_1830 = wire_1672 ^ wire_1671;
assign wire_1831 = wire_1672 & wire_1671;
wire wire_1832, wire_1833;
assign wire_1832 = wire_1674 ^ wire_1673;
assign wire_1833 = wire_1674 & wire_1673;
wire wire_1834, wire_1835;
bit_adder add809(.S(wire_1834), .Cout(wire_1835),  .A(wire_1676), .B(wire_1675), .Cin(wire_1513));
wire wire_1836, wire_1837;
bit_adder add810(.S(wire_1836), .Cout(wire_1837),  .A(wire_1678), .B(wire_1677), .Cin(wire_1515));
wire wire_1838, wire_1839;
bit_adder add811(.S(wire_1838), .Cout(wire_1839),  .A(wire_1680), .B(wire_1679), .Cin(wire_1517));
wire wire_1840, wire_1841;
bit_adder add812(.S(wire_1840), .Cout(wire_1841),  .A(wire_1682), .B(wire_1681), .Cin(wire_1519));
wire wire_1842, wire_1843;
bit_adder add813(.S(wire_1842), .Cout(wire_1843),  .A(wire_1684), .B(wire_1683), .Cin(wire_1521));
wire wire_1844, wire_1845;
bit_adder add814(.S(wire_1844), .Cout(wire_1845),  .A(wire_1686), .B(wire_1685), .Cin(wire_1523));
wire wire_1846, wire_1847;
bit_adder add815(.S(wire_1846), .Cout(wire_1847),  .A(wire_1688), .B(wire_1687), .Cin(wire_1738));
wire wire_1848, wire_1849;
bit_adder add816(.S(wire_1848), .Cout(wire_1849),  .A(wire_1690), .B(wire_1689), .Cin(wire_1740));
wire wire_1850, wire_1851;
bit_adder add817(.S(wire_1850), .Cout(wire_1851),  .A(wire_1692), .B(wire_1691), .Cin(wire_1742));
wire wire_1852, wire_1853;
bit_adder add818(.S(wire_1852), .Cout(wire_1853),  .A(wire_1694), .B(wire_1693), .Cin(wire_1744));
wire wire_1854, wire_1855;
bit_adder add819(.S(wire_1854), .Cout(wire_1855),  .A(wire_1696), .B(wire_1695), .Cin(wire_1746));
wire wire_1856, wire_1857;
bit_adder add820(.S(wire_1856), .Cout(wire_1857),  .A(wire_1698), .B(wire_1697), .Cin(wire_1748));
wire wire_1858, wire_1859;
bit_adder add821(.S(wire_1858), .Cout(wire_1859),  .A(wire_1700), .B(wire_1699), .Cin(wire_1750));
wire wire_1860, wire_1861;
bit_adder add822(.S(wire_1860), .Cout(wire_1861),  .A(wire_1702), .B(wire_1701), .Cin(wire_1752));
wire wire_1862, wire_1863;
bit_adder add823(.S(wire_1862), .Cout(wire_1863),  .A(wire_1704), .B(wire_1703), .Cin(wire_1754));
wire wire_1864, wire_1865;
bit_adder add824(.S(wire_1864), .Cout(wire_1865),  .A(wire_1706), .B(wire_1705), .Cin(wire_1756));
wire wire_1866, wire_1867;
bit_adder add825(.S(wire_1866), .Cout(wire_1867),  .A(wire_1708), .B(wire_1707), .Cin(wire_1758));
wire wire_1868, wire_1869;
bit_adder add826(.S(wire_1868), .Cout(wire_1869),  .A(wire_1710), .B(wire_1709), .Cin(wire_1760));
wire wire_1870, wire_1871;
bit_adder add827(.S(wire_1870), .Cout(wire_1871),  .A(wire_1712), .B(wire_1711), .Cin(wire_1762));
wire wire_1872, wire_1873;
bit_adder add828(.S(wire_1872), .Cout(wire_1873),  .A(wire_1714), .B(wire_1713), .Cin(wire_1764));
wire wire_1874, wire_1875;
bit_adder add829(.S(wire_1874), .Cout(wire_1875),  .A(wire_1716), .B(wire_1715), .Cin(wire_1766));
wire wire_1876, wire_1877;
bit_adder add830(.S(wire_1876), .Cout(wire_1877),  .A(wire_1718), .B(wire_1717), .Cin(wire_1768));
wire wire_1878, wire_1879;
bit_adder add831(.S(wire_1878), .Cout(wire_1879),  .A(wire_1720), .B(wire_1719), .Cin(wire_1770));
wire wire_1880, wire_1881;
bit_adder add832(.S(wire_1880), .Cout(wire_1881),  .A(wire_1722), .B(wire_1721), .Cin(wire_1772));
wire wire_1882, wire_1883;
bit_adder add833(.S(wire_1882), .Cout(wire_1883),  .A(wire_1724), .B(wire_1723), .Cin(wire_1774));
wire wire_1884, wire_1885;
bit_adder add834(.S(wire_1884), .Cout(wire_1885),  .A(wire_1726), .B(wire_1725), .Cin(wire_1776));
wire wire_1886, wire_1887;
bit_adder add835(.S(wire_1886), .Cout(wire_1887),  .A(wire_1728), .B(wire_1727), .Cin(wire_1778));
wire wire_1888, wire_1889;
bit_adder add836(.S(wire_1888), .Cout(wire_1889),  .A(wire_1730), .B(wire_1729), .Cin(wire_1780));
wire wire_1890, wire_1891;
bit_adder add837(.S(wire_1890), .Cout(wire_1891),  .A(wire_1732), .B(wire_1731), .Cin(wire_1782));
wire wire_1892, wire_1893;
bit_adder add838(.S(wire_1892), .Cout(wire_1893),  .A(wire_1734), .B(wire_1733), .Cin(wire_1784));
wire wire_1894, wire_1895;
bit_adder add839(.S(wire_1894), .Cout(wire_1895),  .A(wire_1736), .B(wire_1735), .Cin(wire_1786));
wire wire_1896, wire_1897;
bit_adder add840(.S(wire_1896), .Cout(wire_1897),  .A(wire_1576), .B(wire_1737), .Cin(wire_1788));
wire wire_1898, wire_1899;
assign wire_1898 = wire_1578 ^ wire_1790;
assign wire_1899 = wire_1578 & wire_1790;
wire wire_1900, wire_1901;
assign wire_1900 = wire_1580 ^ wire_1792;
assign wire_1901 = wire_1580 & wire_1792;
wire wire_1902, wire_1903;
assign wire_1902 = wire_1582 ^ wire_1794;
assign wire_1903 = wire_1582 & wire_1794;
wire wire_1904, wire_1905;
assign wire_1904 = wire_1584 ^ wire_1796;
assign wire_1905 = wire_1584 & wire_1796;
wire wire_1906, wire_1907;
assign wire_1906 = wire_966 ^ wire_1798;
assign wire_1907 = wire_966 & wire_1798;
wire wire_1908, wire_1909;
assign wire_1908 = wire_508 ^ wire_1800;
assign wire_1909 = wire_508 & wire_1800;
wire wire_1910, wire_1911;
assign wire_1910 = wire_510 ^ wire_1802;
assign wire_1911 = wire_510 & wire_1802;
wire wire_1912, wire_1913;
assign wire_1912 = partialProduct_23[31] ^ wire_1804;
assign wire_1913 = partialProduct_23[31] & wire_1804;
wire wire_1914, wire_1915;
assign wire_1914 = wire_1818 ^ wire_1817;
assign wire_1915 = wire_1818 & wire_1817;
wire wire_1916, wire_1917;
assign wire_1916 = wire_1820 ^ wire_1819;
assign wire_1917 = wire_1820 & wire_1819;
wire wire_1918, wire_1919;
assign wire_1918 = wire_1822 ^ wire_1821;
assign wire_1919 = wire_1822 & wire_1821;
wire wire_1920, wire_1921;
assign wire_1920 = wire_1824 ^ wire_1823;
assign wire_1921 = wire_1824 & wire_1823;
wire wire_1922, wire_1923;
assign wire_1922 = wire_1826 ^ wire_1825;
assign wire_1923 = wire_1826 & wire_1825;
wire wire_1924, wire_1925;
assign wire_1924 = wire_1828 ^ wire_1827;
assign wire_1925 = wire_1828 & wire_1827;
wire wire_1926, wire_1927;
assign wire_1926 = wire_1830 ^ wire_1829;
assign wire_1927 = wire_1830 & wire_1829;
wire wire_1928, wire_1929;
assign wire_1928 = wire_1832 ^ wire_1831;
assign wire_1929 = wire_1832 & wire_1831;
wire wire_1930, wire_1931;
assign wire_1930 = wire_1834 ^ wire_1833;
assign wire_1931 = wire_1834 & wire_1833;
wire wire_1932, wire_1933;
assign wire_1932 = wire_1836 ^ wire_1835;
assign wire_1933 = wire_1836 & wire_1835;
wire wire_1934, wire_1935;
assign wire_1934 = wire_1838 ^ wire_1837;
assign wire_1935 = wire_1838 & wire_1837;
wire wire_1936, wire_1937;
assign wire_1936 = wire_1840 ^ wire_1839;
assign wire_1937 = wire_1840 & wire_1839;
wire wire_1938, wire_1939;
assign wire_1938 = wire_1842 ^ wire_1841;
assign wire_1939 = wire_1842 & wire_1841;
wire wire_1940, wire_1941;
assign wire_1940 = wire_1844 ^ wire_1843;
assign wire_1941 = wire_1844 & wire_1843;
wire wire_1942, wire_1943;
assign wire_1942 = wire_1846 ^ wire_1845;
assign wire_1943 = wire_1846 & wire_1845;
wire wire_1944, wire_1945;
bit_adder add841(.S(wire_1944), .Cout(wire_1945),  .A(wire_1848), .B(wire_1847), .Cin(wire_1739));
wire wire_1946, wire_1947;
bit_adder add842(.S(wire_1946), .Cout(wire_1947),  .A(wire_1850), .B(wire_1849), .Cin(wire_1741));
wire wire_1948, wire_1949;
bit_adder add843(.S(wire_1948), .Cout(wire_1949),  .A(wire_1852), .B(wire_1851), .Cin(wire_1743));
wire wire_1950, wire_1951;
bit_adder add844(.S(wire_1950), .Cout(wire_1951),  .A(wire_1854), .B(wire_1853), .Cin(wire_1745));
wire wire_1952, wire_1953;
bit_adder add845(.S(wire_1952), .Cout(wire_1953),  .A(wire_1856), .B(wire_1855), .Cin(wire_1747));
wire wire_1954, wire_1955;
bit_adder add846(.S(wire_1954), .Cout(wire_1955),  .A(wire_1858), .B(wire_1857), .Cin(wire_1749));
wire wire_1956, wire_1957;
bit_adder add847(.S(wire_1956), .Cout(wire_1957),  .A(wire_1860), .B(wire_1859), .Cin(wire_1751));
wire wire_1958, wire_1959;
bit_adder add848(.S(wire_1958), .Cout(wire_1959),  .A(wire_1862), .B(wire_1861), .Cin(wire_1753));
wire wire_1960, wire_1961;
bit_adder add849(.S(wire_1960), .Cout(wire_1961),  .A(wire_1864), .B(wire_1863), .Cin(wire_1755));
wire wire_1962, wire_1963;
bit_adder add850(.S(wire_1962), .Cout(wire_1963),  .A(wire_1866), .B(wire_1865), .Cin(wire_1757));
wire wire_1964, wire_1965;
bit_adder add851(.S(wire_1964), .Cout(wire_1965),  .A(wire_1868), .B(wire_1867), .Cin(wire_1759));
wire wire_1966, wire_1967;
bit_adder add852(.S(wire_1966), .Cout(wire_1967),  .A(wire_1870), .B(wire_1869), .Cin(wire_1761));
wire wire_1968, wire_1969;
bit_adder add853(.S(wire_1968), .Cout(wire_1969),  .A(wire_1872), .B(wire_1871), .Cin(wire_1763));
wire wire_1970, wire_1971;
bit_adder add854(.S(wire_1970), .Cout(wire_1971),  .A(wire_1874), .B(wire_1873), .Cin(wire_1765));
wire wire_1972, wire_1973;
bit_adder add855(.S(wire_1972), .Cout(wire_1973),  .A(wire_1876), .B(wire_1875), .Cin(wire_1767));
wire wire_1974, wire_1975;
bit_adder add856(.S(wire_1974), .Cout(wire_1975),  .A(wire_1878), .B(wire_1877), .Cin(wire_1769));
wire wire_1976, wire_1977;
bit_adder add857(.S(wire_1976), .Cout(wire_1977),  .A(wire_1880), .B(wire_1879), .Cin(wire_1771));
wire wire_1978, wire_1979;
bit_adder add858(.S(wire_1978), .Cout(wire_1979),  .A(wire_1882), .B(wire_1881), .Cin(wire_1773));
wire wire_1980, wire_1981;
bit_adder add859(.S(wire_1980), .Cout(wire_1981),  .A(wire_1884), .B(wire_1883), .Cin(wire_1775));
wire wire_1982, wire_1983;
bit_adder add860(.S(wire_1982), .Cout(wire_1983),  .A(wire_1886), .B(wire_1885), .Cin(wire_1777));
wire wire_1984, wire_1985;
bit_adder add861(.S(wire_1984), .Cout(wire_1985),  .A(wire_1888), .B(wire_1887), .Cin(wire_1779));
wire wire_1986, wire_1987;
bit_adder add862(.S(wire_1986), .Cout(wire_1987),  .A(wire_1890), .B(wire_1889), .Cin(wire_1781));
wire wire_1988, wire_1989;
bit_adder add863(.S(wire_1988), .Cout(wire_1989),  .A(wire_1892), .B(wire_1891), .Cin(wire_1783));
wire wire_1990, wire_1991;
bit_adder add864(.S(wire_1990), .Cout(wire_1991),  .A(wire_1894), .B(wire_1893), .Cin(wire_1785));
wire wire_1992, wire_1993;
bit_adder add865(.S(wire_1992), .Cout(wire_1993),  .A(wire_1896), .B(wire_1895), .Cin(wire_1787));
wire wire_1994, wire_1995;
bit_adder add866(.S(wire_1994), .Cout(wire_1995),  .A(wire_1898), .B(wire_1897), .Cin(wire_1789));
wire wire_1996, wire_1997;
bit_adder add867(.S(wire_1996), .Cout(wire_1997),  .A(wire_1900), .B(wire_1899), .Cin(wire_1791));
wire wire_1998, wire_1999;
bit_adder add868(.S(wire_1998), .Cout(wire_1999),  .A(wire_1902), .B(wire_1901), .Cin(wire_1793));
wire wire_2000, wire_2001;
bit_adder add869(.S(wire_2000), .Cout(wire_2001),  .A(wire_1904), .B(wire_1903), .Cin(wire_1795));
wire wire_2002, wire_2003;
bit_adder add870(.S(wire_2002), .Cout(wire_2003),  .A(wire_1906), .B(wire_1905), .Cin(wire_1797));
wire wire_2004, wire_2005;
bit_adder add871(.S(wire_2004), .Cout(wire_2005),  .A(wire_1908), .B(wire_1907), .Cin(wire_1799));
wire wire_2006, wire_2007;
bit_adder add872(.S(wire_2006), .Cout(wire_2007),  .A(wire_1910), .B(wire_1909), .Cin(wire_1801));
wire wire_2008, wire_2009;
bit_adder add873(.S(wire_2008), .Cout(wire_2009),  .A(wire_1912), .B(wire_1911), .Cin(wire_1803));
wire wire_2010, wire_2011;
bit_adder add874(.S(wire_2010), .Cout(wire_2011),  .A(wire_1806), .B(wire_1913), .Cin(wire_1805));
wire wire_2012, wire_2013;
assign wire_2012 = wire_1808 ^ wire_1807;
assign wire_2013 = wire_1808 & wire_1807;
wire wire_2014, wire_2015;
assign wire_2014 = wire_1810 ^ wire_1809;
assign wire_2015 = wire_1810 & wire_1809;
wire wire_2016, wire_2017;
assign wire_2016 = wire_1812 ^ wire_1811;
assign wire_2017 = wire_1812 & wire_1811;
wire wire_2018, wire_2019;
assign wire_2018 = wire_1814 ^ wire_1813;
assign wire_2019 = wire_1814 & wire_1813;
wire wire_2020, wire_2021;
assign wire_2020 = wire_1436 ^ wire_1815;
assign wire_2021 = wire_1436 & wire_1815;
wire wire_2022, wire_2023;
assign wire_2022 = wire_1916 ^ wire_1915;
assign wire_2023 = wire_1916 & wire_1915;
wire wire_2024, wire_2025;
assign wire_2024 = wire_1918 ^ wire_1917;
assign wire_2025 = wire_1918 & wire_1917;
wire wire_2026, wire_2027;
assign wire_2026 = wire_1920 ^ wire_1919;
assign wire_2027 = wire_1920 & wire_1919;
wire wire_2028, wire_2029;
assign wire_2028 = wire_1922 ^ wire_1921;
assign wire_2029 = wire_1922 & wire_1921;
wire wire_2030, wire_2031;
assign wire_2030 = wire_1924 ^ wire_1923;
assign wire_2031 = wire_1924 & wire_1923;
wire wire_2032, wire_2033;
assign wire_2032 = wire_1926 ^ wire_1925;
assign wire_2033 = wire_1926 & wire_1925;
wire wire_2034, wire_2035;
assign wire_2034 = wire_1928 ^ wire_1927;
assign wire_2035 = wire_1928 & wire_1927;
wire wire_2036, wire_2037;
assign wire_2036 = wire_1930 ^ wire_1929;
assign wire_2037 = wire_1930 & wire_1929;
wire wire_2038, wire_2039;
assign wire_2038 = wire_1932 ^ wire_1931;
assign wire_2039 = wire_1932 & wire_1931;
wire wire_2040, wire_2041;
assign wire_2040 = wire_1934 ^ wire_1933;
assign wire_2041 = wire_1934 & wire_1933;
wire wire_2042, wire_2043;
assign wire_2042 = wire_1936 ^ wire_1935;
assign wire_2043 = wire_1936 & wire_1935;
wire wire_2044, wire_2045;
assign wire_2044 = wire_1938 ^ wire_1937;
assign wire_2045 = wire_1938 & wire_1937;
wire wire_2046, wire_2047;
assign wire_2046 = wire_1940 ^ wire_1939;
assign wire_2047 = wire_1940 & wire_1939;
wire wire_2048, wire_2049;
assign wire_2048 = wire_1942 ^ wire_1941;
assign wire_2049 = wire_1942 & wire_1941;
wire wire_2050, wire_2051;
assign wire_2050 = wire_1944 ^ wire_1943;
assign wire_2051 = wire_1944 & wire_1943;
wire wire_2052, wire_2053;
assign wire_2052 = wire_1946 ^ wire_1945;
assign wire_2053 = wire_1946 & wire_1945;
wire wire_2054, wire_2055;
assign wire_2054 = wire_1948 ^ wire_1947;
assign wire_2055 = wire_1948 & wire_1947;
wire wire_2056, wire_2057;
assign wire_2056 = wire_1950 ^ wire_1949;
assign wire_2057 = wire_1950 & wire_1949;
wire wire_2058, wire_2059;
assign wire_2058 = wire_1952 ^ wire_1951;
assign wire_2059 = wire_1952 & wire_1951;
wire wire_2060, wire_2061;
assign wire_2060 = wire_1954 ^ wire_1953;
assign wire_2061 = wire_1954 & wire_1953;
wire wire_2062, wire_2063;
assign wire_2062 = wire_1956 ^ wire_1955;
assign wire_2063 = wire_1956 & wire_1955;
wire wire_2064, wire_2065;
assign wire_2064 = wire_1958 ^ wire_1957;
assign wire_2065 = wire_1958 & wire_1957;
wire wire_2066, wire_2067;
assign wire_2066 = wire_1960 ^ wire_1959;
assign wire_2067 = wire_1960 & wire_1959;
wire wire_2068, wire_2069;
bit_adder add875(.S(wire_2068), .Cout(wire_2069),  .A(wire_1962), .B(wire_1961), .Cin(wire_1377));
wire wire_2070, wire_2071;
bit_adder add876(.S(wire_2070), .Cout(wire_2071),  .A(wire_1964), .B(wire_1963), .Cin(wire_1379));
wire wire_2072, wire_2073;
bit_adder add877(.S(wire_2072), .Cout(wire_2073),  .A(wire_1966), .B(wire_1965), .Cin(wire_1381));
wire wire_2074, wire_2075;
bit_adder add878(.S(wire_2074), .Cout(wire_2075),  .A(wire_1968), .B(wire_1967), .Cin(wire_1383));
wire wire_2076, wire_2077;
bit_adder add879(.S(wire_2076), .Cout(wire_2077),  .A(wire_1970), .B(wire_1969), .Cin(wire_1385));
wire wire_2078, wire_2079;
bit_adder add880(.S(wire_2078), .Cout(wire_2079),  .A(wire_1972), .B(wire_1971), .Cin(wire_1387));
wire wire_2080, wire_2081;
bit_adder add881(.S(wire_2080), .Cout(wire_2081),  .A(wire_1974), .B(wire_1973), .Cin(wire_1389));
wire wire_2082, wire_2083;
bit_adder add882(.S(wire_2082), .Cout(wire_2083),  .A(wire_1976), .B(wire_1975), .Cin(wire_1391));
wire wire_2084, wire_2085;
bit_adder add883(.S(wire_2084), .Cout(wire_2085),  .A(wire_1978), .B(wire_1977), .Cin(wire_1393));
wire wire_2086, wire_2087;
bit_adder add884(.S(wire_2086), .Cout(wire_2087),  .A(wire_1980), .B(wire_1979), .Cin(wire_1395));
wire wire_2088, wire_2089;
bit_adder add885(.S(wire_2088), .Cout(wire_2089),  .A(wire_1982), .B(wire_1981), .Cin(wire_1397));
wire wire_2090, wire_2091;
bit_adder add886(.S(wire_2090), .Cout(wire_2091),  .A(wire_1984), .B(wire_1983), .Cin(wire_1399));
wire wire_2092, wire_2093;
bit_adder add887(.S(wire_2092), .Cout(wire_2093),  .A(wire_1986), .B(wire_1985), .Cin(wire_1401));
wire wire_2094, wire_2095;
bit_adder add888(.S(wire_2094), .Cout(wire_2095),  .A(wire_1988), .B(wire_1987), .Cin(wire_1403));
wire wire_2096, wire_2097;
bit_adder add889(.S(wire_2096), .Cout(wire_2097),  .A(wire_1990), .B(wire_1989), .Cin(wire_1405));
wire wire_2098, wire_2099;
bit_adder add890(.S(wire_2098), .Cout(wire_2099),  .A(wire_1992), .B(wire_1991), .Cin(wire_1407));
wire wire_2100, wire_2101;
bit_adder add891(.S(wire_2100), .Cout(wire_2101),  .A(wire_1994), .B(wire_1993), .Cin(wire_1409));
wire wire_2102, wire_2103;
bit_adder add892(.S(wire_2102), .Cout(wire_2103),  .A(wire_1996), .B(wire_1995), .Cin(wire_1411));
wire wire_2104, wire_2105;
bit_adder add893(.S(wire_2104), .Cout(wire_2105),  .A(wire_1998), .B(wire_1997), .Cin(wire_1413));
wire wire_2106, wire_2107;
bit_adder add894(.S(wire_2106), .Cout(wire_2107),  .A(wire_2000), .B(wire_1999), .Cin(wire_1415));
wire wire_2108, wire_2109;
bit_adder add895(.S(wire_2108), .Cout(wire_2109),  .A(wire_2002), .B(wire_2001), .Cin(wire_1417));
wire wire_2110, wire_2111;
bit_adder add896(.S(wire_2110), .Cout(wire_2111),  .A(wire_2004), .B(wire_2003), .Cin(wire_1419));
wire wire_2112, wire_2113;
bit_adder add897(.S(wire_2112), .Cout(wire_2113),  .A(wire_2006), .B(wire_2005), .Cin(wire_1421));
wire wire_2114, wire_2115;
bit_adder add898(.S(wire_2114), .Cout(wire_2115),  .A(wire_2008), .B(wire_2007), .Cin(wire_1423));
wire wire_2116, wire_2117;
bit_adder add899(.S(wire_2116), .Cout(wire_2117),  .A(wire_2010), .B(wire_2009), .Cin(wire_1425));
wire wire_2118, wire_2119;
bit_adder add900(.S(wire_2118), .Cout(wire_2119),  .A(wire_2012), .B(wire_2011), .Cin(wire_1427));
wire wire_2120, wire_2121;
bit_adder add901(.S(wire_2120), .Cout(wire_2121),  .A(wire_2014), .B(wire_2013), .Cin(wire_1429));
wire wire_2122, wire_2123;
bit_adder add902(.S(wire_2122), .Cout(wire_2123),  .A(wire_2016), .B(wire_2015), .Cin(wire_1431));
wire wire_2124, wire_2125;
bit_adder add903(.S(wire_2124), .Cout(wire_2125),  .A(wire_2018), .B(wire_2017), .Cin(wire_1433));
wire wire_2126, wire_2127;
bit_adder add904(.S(wire_2126), .Cout(wire_2127),  .A(wire_2020), .B(wire_2019), .Cin(wire_1435));
wire wire_2128, wire_2129;
bit_adder add905(.S(wire_2128), .Cout(wire_2129),  .A(wire_1438), .B(wire_2021), .Cin(wire_1437));
wire wire_2130, wire_2131;
assign wire_2130 = partialProduct_31[31] ^ wire_1439;
assign wire_2131 = partialProduct_31[31] & wire_1439;
// Final combination
wire wire_2132, wire_2133;
bit_adder add906(.S(wire_2132), .Cout(wire_2133),  .A(wire_2024), .B(wire_2023), .Cin(1'b0));
wire wire_2134, wire_2135;
bit_adder add907(.S(wire_2134), .Cout(wire_2135),  .A(wire_2026), .B(wire_2025), .Cin(wire_2133));
wire wire_2136, wire_2137;
bit_adder add908(.S(wire_2136), .Cout(wire_2137),  .A(wire_2028), .B(wire_2027), .Cin(wire_2135));
wire wire_2138, wire_2139;
bit_adder add909(.S(wire_2138), .Cout(wire_2139),  .A(wire_2030), .B(wire_2029), .Cin(wire_2137));
wire wire_2140, wire_2141;
bit_adder add910(.S(wire_2140), .Cout(wire_2141),  .A(wire_2032), .B(wire_2031), .Cin(wire_2139));
wire wire_2142, wire_2143;
bit_adder add911(.S(wire_2142), .Cout(wire_2143),  .A(wire_2034), .B(wire_2033), .Cin(wire_2141));
wire wire_2144, wire_2145;
bit_adder add912(.S(wire_2144), .Cout(wire_2145),  .A(wire_2036), .B(wire_2035), .Cin(wire_2143));
wire wire_2146, wire_2147;
bit_adder add913(.S(wire_2146), .Cout(wire_2147),  .A(wire_2038), .B(wire_2037), .Cin(wire_2145));
wire wire_2148, wire_2149;
bit_adder add914(.S(wire_2148), .Cout(wire_2149),  .A(wire_2040), .B(wire_2039), .Cin(wire_2147));
wire wire_2150, wire_2151;
bit_adder add915(.S(wire_2150), .Cout(wire_2151),  .A(wire_2042), .B(wire_2041), .Cin(wire_2149));
wire wire_2152, wire_2153;
bit_adder add916(.S(wire_2152), .Cout(wire_2153),  .A(wire_2044), .B(wire_2043), .Cin(wire_2151));
wire wire_2154, wire_2155;
bit_adder add917(.S(wire_2154), .Cout(wire_2155),  .A(wire_2046), .B(wire_2045), .Cin(wire_2153));
wire wire_2156, wire_2157;
bit_adder add918(.S(wire_2156), .Cout(wire_2157),  .A(wire_2048), .B(wire_2047), .Cin(wire_2155));
wire wire_2158, wire_2159;
bit_adder add919(.S(wire_2158), .Cout(wire_2159),  .A(wire_2050), .B(wire_2049), .Cin(wire_2157));
wire wire_2160, wire_2161;
bit_adder add920(.S(wire_2160), .Cout(wire_2161),  .A(wire_2052), .B(wire_2051), .Cin(wire_2159));
wire wire_2162, wire_2163;
bit_adder add921(.S(wire_2162), .Cout(wire_2163),  .A(wire_2054), .B(wire_2053), .Cin(wire_2161));
wire wire_2164, wire_2165;
bit_adder add922(.S(wire_2164), .Cout(wire_2165),  .A(wire_2056), .B(wire_2055), .Cin(wire_2163));
wire wire_2166, wire_2167;
bit_adder add923(.S(wire_2166), .Cout(wire_2167),  .A(wire_2058), .B(wire_2057), .Cin(wire_2165));
wire wire_2168, wire_2169;
bit_adder add924(.S(wire_2168), .Cout(wire_2169),  .A(wire_2060), .B(wire_2059), .Cin(wire_2167));
wire wire_2170, wire_2171;
bit_adder add925(.S(wire_2170), .Cout(wire_2171),  .A(wire_2062), .B(wire_2061), .Cin(wire_2169));
wire wire_2172, wire_2173;
bit_adder add926(.S(wire_2172), .Cout(wire_2173),  .A(wire_2064), .B(wire_2063), .Cin(wire_2171));
wire wire_2174, wire_2175;
bit_adder add927(.S(wire_2174), .Cout(wire_2175),  .A(wire_2066), .B(wire_2065), .Cin(wire_2173));
wire wire_2176, wire_2177;
bit_adder add928(.S(wire_2176), .Cout(wire_2177),  .A(wire_2068), .B(wire_2067), .Cin(wire_2175));
wire wire_2178, wire_2179;
bit_adder add929(.S(wire_2178), .Cout(wire_2179),  .A(wire_2070), .B(wire_2069), .Cin(wire_2177));
wire wire_2180, wire_2181;
bit_adder add930(.S(wire_2180), .Cout(wire_2181),  .A(wire_2072), .B(wire_2071), .Cin(wire_2179));
wire wire_2182, wire_2183;
bit_adder add931(.S(wire_2182), .Cout(wire_2183),  .A(wire_2074), .B(wire_2073), .Cin(wire_2181));
wire wire_2184, wire_2185;
bit_adder add932(.S(wire_2184), .Cout(wire_2185),  .A(wire_2076), .B(wire_2075), .Cin(wire_2183));
wire wire_2186, wire_2187;
bit_adder add933(.S(wire_2186), .Cout(wire_2187),  .A(wire_2078), .B(wire_2077), .Cin(wire_2185));
wire wire_2188, wire_2189;
bit_adder add934(.S(wire_2188), .Cout(wire_2189),  .A(wire_2080), .B(wire_2079), .Cin(wire_2187));
wire wire_2190, wire_2191;
bit_adder add935(.S(wire_2190), .Cout(wire_2191),  .A(wire_2082), .B(wire_2081), .Cin(wire_2189));
wire wire_2192, wire_2193;
bit_adder add936(.S(wire_2192), .Cout(wire_2193),  .A(wire_2084), .B(wire_2083), .Cin(wire_2191));
wire wire_2194, wire_2195;
bit_adder add937(.S(wire_2194), .Cout(wire_2195),  .A(wire_2086), .B(wire_2085), .Cin(wire_2193));
wire wire_2196, wire_2197;
bit_adder add938(.S(wire_2196), .Cout(wire_2197),  .A(wire_2088), .B(wire_2087), .Cin(wire_2195));
wire wire_2198, wire_2199;
bit_adder add939(.S(wire_2198), .Cout(wire_2199),  .A(wire_2090), .B(wire_2089), .Cin(wire_2197));
wire wire_2200, wire_2201;
bit_adder add940(.S(wire_2200), .Cout(wire_2201),  .A(wire_2092), .B(wire_2091), .Cin(wire_2199));
wire wire_2202, wire_2203;
bit_adder add941(.S(wire_2202), .Cout(wire_2203),  .A(wire_2094), .B(wire_2093), .Cin(wire_2201));
wire wire_2204, wire_2205;
bit_adder add942(.S(wire_2204), .Cout(wire_2205),  .A(wire_2096), .B(wire_2095), .Cin(wire_2203));
wire wire_2206, wire_2207;
bit_adder add943(.S(wire_2206), .Cout(wire_2207),  .A(wire_2098), .B(wire_2097), .Cin(wire_2205));
wire wire_2208, wire_2209;
bit_adder add944(.S(wire_2208), .Cout(wire_2209),  .A(wire_2100), .B(wire_2099), .Cin(wire_2207));
wire wire_2210, wire_2211;
bit_adder add945(.S(wire_2210), .Cout(wire_2211),  .A(wire_2102), .B(wire_2101), .Cin(wire_2209));
wire wire_2212, wire_2213;
bit_adder add946(.S(wire_2212), .Cout(wire_2213),  .A(wire_2104), .B(wire_2103), .Cin(wire_2211));
wire wire_2214, wire_2215;
bit_adder add947(.S(wire_2214), .Cout(wire_2215),  .A(wire_2106), .B(wire_2105), .Cin(wire_2213));
wire wire_2216, wire_2217;
bit_adder add948(.S(wire_2216), .Cout(wire_2217),  .A(wire_2108), .B(wire_2107), .Cin(wire_2215));
wire wire_2218, wire_2219;
bit_adder add949(.S(wire_2218), .Cout(wire_2219),  .A(wire_2110), .B(wire_2109), .Cin(wire_2217));
wire wire_2220, wire_2221;
bit_adder add950(.S(wire_2220), .Cout(wire_2221),  .A(wire_2112), .B(wire_2111), .Cin(wire_2219));
wire wire_2222, wire_2223;
bit_adder add951(.S(wire_2222), .Cout(wire_2223),  .A(wire_2114), .B(wire_2113), .Cin(wire_2221));
wire wire_2224, wire_2225;
bit_adder add952(.S(wire_2224), .Cout(wire_2225),  .A(wire_2116), .B(wire_2115), .Cin(wire_2223));
wire wire_2226, wire_2227;
bit_adder add953(.S(wire_2226), .Cout(wire_2227),  .A(wire_2118), .B(wire_2117), .Cin(wire_2225));
wire wire_2228, wire_2229;
bit_adder add954(.S(wire_2228), .Cout(wire_2229),  .A(wire_2120), .B(wire_2119), .Cin(wire_2227));
wire wire_2230, wire_2231;
bit_adder add955(.S(wire_2230), .Cout(wire_2231),  .A(wire_2122), .B(wire_2121), .Cin(wire_2229));
wire wire_2232, wire_2233;
bit_adder add956(.S(wire_2232), .Cout(wire_2233),  .A(wire_2124), .B(wire_2123), .Cin(wire_2231));
wire wire_2234, wire_2235;
bit_adder add957(.S(wire_2234), .Cout(wire_2235),  .A(wire_2126), .B(wire_2125), .Cin(wire_2233));
wire wire_2236, wire_2237;
bit_adder add958(.S(wire_2236), .Cout(wire_2237),  .A(wire_2128), .B(wire_2127), .Cin(wire_2235));
wire wire_2238, wire_2239;
bit_adder add959(.S(wire_2238), .Cout(wire_2239),  .A(wire_2130), .B(wire_2129), .Cin(wire_2237));
assign data_result[0] = partialProduct_0[0];
assign data_result[1] = wire_0;
assign data_result[2] = wire_640;
assign data_result[3] = wire_1100;
assign data_result[4] = wire_1440;
assign data_result[5] = wire_1656;
assign data_result[6] = wire_1816;
assign data_result[7] = wire_1914;
assign data_result[8] = wire_2022;
assign data_result[9] = wire_2132;
assign data_result[10] = wire_2134;
assign data_result[11] = wire_2136;
assign data_result[12] = wire_2138;
assign data_result[13] = wire_2140;
assign data_result[14] = wire_2142;
assign data_result[15] = wire_2144;
assign data_result[16] = wire_2146;
assign data_result[17] = wire_2148;
assign data_result[18] = wire_2150;
assign data_result[19] = wire_2152;
assign data_result[20] = wire_2154;
assign data_result[21] = wire_2156;
assign data_result[22] = wire_2158;
assign data_result[23] = wire_2160;
assign data_result[24] = wire_2162;
assign data_result[25] = wire_2164;
assign data_result[26] = wire_2166;
assign data_result[27] = wire_2168;
assign data_result[28] = wire_2170;
assign data_result[29] = wire_2172;
assign data_result[30] = wire_2174;
assign data_result[31] = wire_2176;
assign data_result[32] = wire_2178;
assign data_result[33] = wire_2180;
assign data_result[34] = wire_2182;
assign data_result[35] = wire_2184;
assign data_result[36] = wire_2186;
assign data_result[37] = wire_2188;
assign data_result[38] = wire_2190;
assign data_result[39] = wire_2192;
assign data_result[40] = wire_2194;
assign data_result[41] = wire_2196;
assign data_result[42] = wire_2198;
assign data_result[43] = wire_2200;
assign data_result[44] = wire_2202;
assign data_result[45] = wire_2204;
assign data_result[46] = wire_2206;
assign data_result[47] = wire_2208;
assign data_result[48] = wire_2210;
assign data_result[49] = wire_2212;
assign data_result[50] = wire_2214;
assign data_result[51] = wire_2216;
assign data_result[52] = wire_2218;
assign data_result[53] = wire_2220;
assign data_result[54] = wire_2222;
assign data_result[55] = wire_2224;
assign data_result[56] = wire_2226;
assign data_result[57] = wire_2228;
assign data_result[58] = wire_2230;
assign data_result[59] = wire_2232;
assign data_result[60] = wire_2234;
assign data_result[61] = wire_2236;
assign data_result[62] = wire_2238;
wire burner;
assign data_result[63] = wire_2239;

wire andOverflow, orOverflow;
assign andOverflow = &data_result[63:31];
assign orOverflow = |data_result[63:31];
assign data_exception = (!andOverflow) & (orOverflow);

endmodule
