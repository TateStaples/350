module decode32(out, ctrl)
    input [4:0] ctrl;
    output [31:0] out;

    

    and and0(out[0], );
endmodule