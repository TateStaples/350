module divider(
    data_operandA, data_operandB, // inputs
    clock, ctrl_DIV, // control
    data_quotient, data_remainder, data_exception, data_resultRDY);  // outputs

endmodule